----------------------------------------------------------------------------------
-- Company: ECL - Institut des Nanotechnologies de Lyon
-- Engineer: MATRANGOLO Paul-Antoine
-- 
-- Create Date: 09.03.2021 15:46:44
-- Design Name: FeFET Emulator
-- Module Name: tb_FeFET_nand - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: This testbench aim to test de FeFET component to get output tension
-- and behavioral simulation.
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE; use IEEE.STD_LOGIC_1164.ALL;
-- Uncomment the following library declaration if using 
-- arithmetic functions with Signed or Unsigned values 
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating 
-- any Xilinx leaf cells in this code. 
--library UNISIM; 
--use UNISIM.VComponents.all;

library ieee_proposed;
use ieee_proposed.fixed_float_types.all;
use ieee_proposed.fixed_pkg.all;

entity Simul1 is 
-- Port ( ); 
end Simul1;

architecture Behavioral of Simul1 is
    component FeFET1 is 
        Port (  Vi : in std_logic_vector(23 downto 0);
                Vo : out std_logic_vector(23 downto 0));
    end component FeFET1;
    
    signal Vin : std_logic_vector(23 downto 0) := X"000000"; 
    signal Vout : std_logic_vector(23 downto 0);
     
begin
    FF1 : FeFET1 port map ( Vi => Vin, Vo => Vout);
    
    -- this testbench was generated with a function in Python

    -- double ramp
    Vin <= X"800000" after 0.0us,
    X"808312" after 0.2002002002002002us,
    X"810624" after 0.4004004004004004us,
    X"818937" after 0.6006006006006006us,
    X"820c49" after 0.8008008008008008us,
    X"828f5c" after 1.001001001001001us,
    X"83126e" after 1.2012012012012012us,
    X"839580" after 1.4014014014014016us,
    X"841893" after 1.6016016016016017us,
    X"849ba5" after 1.8018018018018018us,
    X"851eb8" after 2.002002002002002us,
    X"85a1ca" after 2.2022022022022023us,
    X"8624dd" after 2.4024024024024024us,
    X"86a7ef" after 2.6026026026026026us,
    X"872b01" after 2.802802802802803us,
    X"87ae14" after 3.0030030030030033us,
    X"883126" after 3.2032032032032034us,
    X"88b439" after 3.4034034034034035us,
    X"89374b" after 3.6036036036036037us,
    X"89ba5e" after 3.8038038038038042us,
    X"8a3d70" after 4.004004004004004us,
    X"8ac082" after 4.2042042042042045us,
    X"8b4395" after 4.404404404404405us,
    X"8bc6a7" after 4.604604604604605us,
    X"8c49ba" after 4.804804804804805us,
    X"8ccccc" after 5.005005005005005us,
    X"8d4fdf" after 5.205205205205205us,
    X"8dd2f1" after 5.405405405405406us,
    X"8e5603" after 5.605605605605606us,
    X"8ed916" after 5.805805805805806us,
    X"8f5c28" after 6.0060060060060065us,
    X"8fdf3b" after 6.206206206206207us,
    X"90624d" after 6.406406406406407us,
    X"90e560" after 6.606606606606607us,
    X"916872" after 6.806806806806807us,
    X"91eb84" after 7.007007007007007us,
    X"926e97" after 7.207207207207207us,
    X"92f1a9" after 7.407407407407407us,
    X"9374bc" after 7.6076076076076085us,
    X"93f7ce" after 7.807807807807809us,
    X"947ae1" after 8.008008008008009us,
    X"94fdf3" after 8.208208208208209us,
    X"958105" after 8.408408408408409us,
    X"960418" after 8.608608608608609us,
    X"96872a" after 8.80880880880881us,
    X"970a3d" after 9.00900900900901us,
    X"978d4f" after 9.20920920920921us,
    X"981062" after 9.40940940940941us,
    X"989374" after 9.60960960960961us,
    X"991686" after 9.80980980980981us,
    X"999999" after 10.01001001001001us,
    X"9a1cab" after 10.21021021021021us,
    X"9a9fbe" after 10.41041041041041us,
    X"9b22d0" after 10.61061061061061us,
    X"9ba5e3" after 10.810810810810812us,
    X"9c28f5" after 11.011011011011012us,
    X"9cac07" after 11.211211211211213us,
    X"9d2f1a" after 11.411411411411413us,
    X"9db22c" after 11.611611611611613us,
    X"9e353f" after 11.811811811811813us,
    X"9eb851" after 12.012012012012013us,
    X"9f3b64" after 12.212212212212213us,
    X"9fbe76" after 12.412412412412413us,
    X"a04188" after 12.612612612612613us,
    X"a0c49b" after 12.812812812812814us,
    X"a147ad" after 13.013013013013014us,
    X"a1cac0" after 13.213213213213214us,
    X"a24dd2" after 13.413413413413414us,
    X"a2d0e5" after 13.613613613613614us,
    X"a353f7" after 13.813813813813814us,
    X"a3d709" after 14.014014014014014us,
    X"a45a1c" after 14.214214214214214us,
    X"a4dd2e" after 14.414414414414415us,
    X"a56041" after 14.614614614614615us,
    X"a5e353" after 14.814814814814815us,
    X"a66666" after 15.015015015015017us,
    X"a6e978" after 15.215215215215217us,
    X"a76c8a" after 15.415415415415417us,
    X"a7ef9d" after 15.615615615615617us,
    X"a872af" after 15.815815815815817us,
    X"a8f5c2" after 16.016016016016017us,
    X"a978d4" after 16.216216216216218us,
    X"a9fbe7" after 16.416416416416418us,
    X"aa7ef9" after 16.616616616616618us,
    X"ab020b" after 16.816816816816818us,
    X"ab851e" after 17.017017017017018us,
    X"ac0830" after 17.217217217217218us,
    X"ac8b43" after 17.41741741741742us,
    X"ad0e55" after 17.61761761761762us,
    X"ad9168" after 17.81781781781782us,
    X"ae147a" after 18.01801801801802us,
    X"ae978c" after 18.21821821821822us,
    X"af1a9f" after 18.41841841841842us,
    X"af9db1" after 18.61861861861862us,
    X"b020c4" after 18.81881881881882us,
    X"b0a3d6" after 19.01901901901902us,
    X"b126e9" after 19.21921921921922us,
    X"b1a9fb" after 19.41941941941942us,
    X"b22d0d" after 19.61961961961962us,
    X"b2b020" after 19.81981981981982us,
    X"b33332" after 20.02002002002002us,
    X"b3b645" after 20.22022022022022us,
    X"b43957" after 20.42042042042042us,
    X"b4bc6a" after 20.62062062062062us,
    X"b53f7c" after 20.82082082082082us,
    X"b5c28e" after 21.02102102102102us,
    X"b645a1" after 21.22122122122122us,
    X"b6c8b3" after 21.421421421421424us,
    X"b74bc6" after 21.621621621621625us,
    X"b7ced8" after 21.821821821821825us,
    X"b851eb" after 22.022022022022025us,
    X"b8d4fd" after 22.222222222222225us,
    X"b9580f" after 22.422422422422425us,
    X"b9db22" after 22.622622622622625us,
    X"ba5e34" after 22.822822822822825us,
    X"bae147" after 23.023023023023026us,
    X"bb6459" after 23.223223223223226us,
    X"bbe76c" after 23.423423423423426us,
    X"bc6a7e" after 23.623623623623626us,
    X"bced90" after 23.823823823823826us,
    X"bd70a3" after 24.024024024024026us,
    X"bdf3b5" after 24.224224224224226us,
    X"be76c8" after 24.424424424424426us,
    X"bef9da" after 24.624624624624627us,
    X"bf7ced" after 24.824824824824827us,
    X"bfffff" after 25.025025025025027us,
    X"c08311" after 25.225225225225227us,
    X"c10624" after 25.425425425425427us,
    X"c18936" after 25.625625625625627us,
    X"c20c49" after 25.825825825825827us,
    X"c28f5b" after 26.026026026026027us,
    X"c3126e" after 26.226226226226228us,
    X"c39580" after 26.426426426426428us,
    X"c41892" after 26.626626626626628us,
    X"c49ba5" after 26.826826826826828us,
    X"c51eb7" after 27.027027027027028us,
    X"c5a1ca" after 27.227227227227228us,
    X"c624dc" after 27.42742742742743us,
    X"c6a7ef" after 27.62762762762763us,
    X"c72b01" after 27.82782782782783us,
    X"c7ae13" after 28.02802802802803us,
    X"c83126" after 28.22822822822823us,
    X"c8b438" after 28.42842842842843us,
    X"c9374b" after 28.62862862862863us,
    X"c9ba5d" after 28.82882882882883us,
    X"ca3d70" after 29.02902902902903us,
    X"cac082" after 29.22922922922923us,
    X"cb4394" after 29.42942942942943us,
    X"cbc6a7" after 29.62962962962963us,
    X"cc49b9" after 29.82982982982983us,
    X"cccccc" after 30.030030030030034us,
    X"cd4fde" after 30.230230230230234us,
    X"cdd2f1" after 30.430430430430434us,
    X"ce5603" after 30.630630630630634us,
    X"ced915" after 30.830830830830834us,
    X"cf5c28" after 31.031031031031034us,
    X"cfdf3a" after 31.231231231231234us,
    X"d0624d" after 31.431431431431434us,
    X"d0e55f" after 31.631631631631635us,
    X"d16872" after 31.831831831831835us,
    X"d1eb84" after 32.032032032032035us,
    X"d26e96" after 32.232232232232235us,
    X"d2f1a9" after 32.432432432432435us,
    X"d374bb" after 32.632632632632635us,
    X"d3f7ce" after 32.832832832832835us,
    X"d47ae0" after 33.033033033033036us,
    X"d4fdf3" after 33.233233233233236us,
    X"d58105" after 33.433433433433436us,
    X"d60417" after 33.633633633633636us,
    X"d6872a" after 33.833833833833836us,
    X"d70a3c" after 34.034034034034036us,
    X"d78d4f" after 34.234234234234236us,
    X"d81061" after 34.434434434434436us,
    X"d89374" after 34.63463463463464us,
    X"d91686" after 34.83483483483484us,
    X"d99998" after 35.03503503503504us,
    X"da1cab" after 35.23523523523524us,
    X"da9fbd" after 35.43543543543544us,
    X"db22d0" after 35.63563563563564us,
    X"dba5e2" after 35.83583583583584us,
    X"dc28f5" after 36.03603603603604us,
    X"dcac07" after 36.23623623623624us,
    X"dd2f19" after 36.43643643643644us,
    X"ddb22c" after 36.63663663663664us,
    X"de353e" after 36.83683683683684us,
    X"deb851" after 37.03703703703704us,
    X"df3b63" after 37.23723723723724us,
    X"dfbe76" after 37.43743743743744us,
    X"e04188" after 37.63763763763764us,
    X"e0c49a" after 37.83783783783784us,
    X"e147ad" after 38.03803803803804us,
    X"e1cabf" after 38.23823823823824us,
    X"e24dd2" after 38.43843843843844us,
    X"e2d0e4" after 38.63863863863864us,
    X"e353f7" after 38.83883883883884us,
    X"e3d709" after 39.03903903903904us,
    X"e45a1b" after 39.23923923923924us,
    X"e4dd2e" after 39.43943943943944us,
    X"e56040" after 39.63963963963964us,
    X"e5e353" after 39.83983983983984us,
    X"e66665" after 40.04004004004004us,
    X"e6e978" after 40.24024024024024us,
    X"e76c8a" after 40.44044044044044us,
    X"e7ef9c" after 40.64064064064064us,
    X"e872af" after 40.84084084084084us,
    X"e8f5c1" after 41.04104104104104us,
    X"e978d4" after 41.24124124124124us,
    X"e9fbe6" after 41.44144144144144us,
    X"ea7ef9" after 41.64164164164164us,
    X"eb020b" after 41.84184184184184us,
    X"eb851d" after 42.04204204204204us,
    X"ec0830" after 42.24224224224224us,
    X"ec8b42" after 42.44244244244244us,
    X"ed0e55" after 42.64264264264264us,
    X"ed9167" after 42.84284284284285us,
    X"ee147a" after 43.04304304304305us,
    X"ee978c" after 43.24324324324325us,
    X"ef1a9e" after 43.44344344344345us,
    X"ef9db1" after 43.64364364364365us,
    X"f020c3" after 43.84384384384385us,
    X"f0a3d6" after 44.04404404404405us,
    X"f126e8" after 44.24424424424425us,
    X"f1a9fb" after 44.44444444444445us,
    X"f22d0d" after 44.64464464464465us,
    X"f2b01f" after 44.84484484484485us,
    X"f33332" after 45.04504504504505us,
    X"f3b644" after 45.24524524524525us,
    X"f43957" after 45.44544544544545us,
    X"f4bc69" after 45.64564564564565us,
    X"f53f7c" after 45.84584584584585us,
    X"f5c28e" after 46.04604604604605us,
    X"f645a0" after 46.24624624624625us,
    X"f6c8b3" after 46.44644644644645us,
    X"f74bc5" after 46.64664664664665us,
    X"f7ced8" after 46.84684684684685us,
    X"f851ea" after 47.04704704704705us,
    X"f8d4fd" after 47.24724724724725us,
    X"f9580f" after 47.44744744744745us,
    X"f9db21" after 47.64764764764765us,
    X"fa5e34" after 47.84784784784785us,
    X"fae146" after 48.04804804804805us,
    X"fb6459" after 48.24824824824825us,
    X"fbe76b" after 48.44844844844845us,
    X"fc6a7e" after 48.64864864864865us,
    X"fced90" after 48.84884884884885us,
    X"fd70a2" after 49.04904904904905us,
    X"fdf3b5" after 49.24924924924925us,
    X"fe76c7" after 49.44944944944945us,
    X"fef9da" after 49.64964964964965us,
    X"ff7cec" after 49.84984984984985us,
    X"000000" after 50.050050050050054us,
    X"008312" after 50.250250250250254us,
    X"010624" after 50.450450450450454us,
    X"018937" after 50.650650650650654us,
    X"020c49" after 50.850850850850854us,
    X"028f5c" after 51.051051051051054us,
    X"03126e" after 51.251251251251254us,
    X"039580" after 51.451451451451454us,
    X"041893" after 51.651651651651655us,
    X"049ba5" after 51.851851851851855us,
    X"051eb8" after 52.052052052052055us,
    X"05a1ca" after 52.252252252252255us,
    X"0624dd" after 52.452452452452455us,
    X"06a7ef" after 52.652652652652655us,
    X"072b01" after 52.852852852852855us,
    X"07ae14" after 53.053053053053056us,
    X"083126" after 53.253253253253256us,
    X"08b439" after 53.453453453453456us,
    X"09374b" after 53.653653653653656us,
    X"09ba5e" after 53.853853853853856us,
    X"0a3d70" after 54.054054054054056us,
    X"0ac082" after 54.254254254254256us,
    X"0b4395" after 54.454454454454456us,
    X"0bc6a7" after 54.65465465465466us,
    X"0c49ba" after 54.85485485485486us,
    X"0ccccc" after 55.05505505505506us,
    X"0d4fdf" after 55.25525525525526us,
    X"0dd2f1" after 55.45545545545546us,
    X"0e5603" after 55.65565565565566us,
    X"0ed916" after 55.85585585585586us,
    X"0f5c28" after 56.05605605605606us,
    X"0fdf3b" after 56.25625625625626us,
    X"10624d" after 56.45645645645646us,
    X"10e560" after 56.65665665665666us,
    X"116872" after 56.85685685685686us,
    X"11eb84" after 57.05705705705706us,
    X"126e97" after 57.25725725725726us,
    X"12f1a9" after 57.45745745745746us,
    X"1374bc" after 57.65765765765766us,
    X"13f7ce" after 57.85785785785786us,
    X"147ae1" after 58.05805805805806us,
    X"14fdf3" after 58.25825825825826us,
    X"158105" after 58.45845845845846us,
    X"160418" after 58.65865865865866us,
    X"16872a" after 58.85885885885886us,
    X"170a3d" after 59.05905905905906us,
    X"178d4f" after 59.25925925925926us,
    X"181062" after 59.45945945945946us,
    X"189374" after 59.65965965965966us,
    X"191686" after 59.85985985985987us,
    X"199999" after 60.06006006006007us,
    X"1a1cab" after 60.26026026026027us,
    X"1a9fbe" after 60.46046046046047us,
    X"1b22d0" after 60.66066066066067us,
    X"1ba5e3" after 60.86086086086087us,
    X"1c28f5" after 61.06106106106107us,
    X"1cac07" after 61.26126126126127us,
    X"1d2f1a" after 61.46146146146147us,
    X"1db22c" after 61.66166166166167us,
    X"1e353f" after 61.86186186186187us,
    X"1eb851" after 62.06206206206207us,
    X"1f3b64" after 62.26226226226227us,
    X"1fbe76" after 62.46246246246247us,
    X"204188" after 62.66266266266267us,
    X"20c49b" after 62.86286286286287us,
    X"2147ad" after 63.06306306306307us,
    X"21cac0" after 63.26326326326327us,
    X"224dd2" after 63.46346346346347us,
    X"22d0e5" after 63.66366366366367us,
    X"2353f7" after 63.86386386386387us,
    X"23d709" after 64.06406406406407us,
    X"245a1c" after 64.26426426426427us,
    X"24dd2e" after 64.46446446446447us,
    X"256041" after 64.66466466466467us,
    X"25e353" after 64.86486486486487us,
    X"266666" after 65.06506506506507us,
    X"26e978" after 65.26526526526527us,
    X"276c8a" after 65.46546546546547us,
    X"27ef9d" after 65.66566566566567us,
    X"2872af" after 65.86586586586587us,
    X"28f5c2" after 66.06606606606607us,
    X"2978d4" after 66.26626626626627us,
    X"29fbe7" after 66.46646646646647us,
    X"2a7ef9" after 66.66666666666667us,
    X"2b020b" after 66.86686686686687us,
    X"2b851e" after 67.06706706706707us,
    X"2c0830" after 67.26726726726727us,
    X"2c8b43" after 67.46746746746747us,
    X"2d0e55" after 67.66766766766767us,
    X"2d9168" after 67.86786786786787us,
    X"2e147a" after 68.06806806806807us,
    X"2e978c" after 68.26826826826827us,
    X"2f1a9f" after 68.46846846846847us,
    X"2f9db1" after 68.66866866866867us,
    X"3020c4" after 68.86886886886887us,
    X"30a3d6" after 69.06906906906907us,
    X"3126e9" after 69.26926926926927us,
    X"31a9fb" after 69.46946946946947us,
    X"322d0d" after 69.66966966966967us,
    X"32b020" after 69.86986986986987us,
    X"333332" after 70.07007007007007us,
    X"33b645" after 70.27027027027027us,
    X"343957" after 70.47047047047047us,
    X"34bc6a" after 70.67067067067067us,
    X"353f7c" after 70.87087087087087us,
    X"35c28e" after 71.07107107107107us,
    X"3645a1" after 71.27127127127127us,
    X"36c8b3" after 71.47147147147147us,
    X"374bc6" after 71.67167167167167us,
    X"37ced8" after 71.87187187187187us,
    X"3851eb" after 72.07207207207207us,
    X"38d4fd" after 72.27227227227228us,
    X"39580f" after 72.47247247247248us,
    X"39db22" after 72.67267267267268us,
    X"3a5e34" after 72.87287287287288us,
    X"3ae147" after 73.07307307307308us,
    X"3b6459" after 73.27327327327328us,
    X"3be76c" after 73.47347347347348us,
    X"3c6a7e" after 73.67367367367368us,
    X"3ced90" after 73.87387387387388us,
    X"3d70a3" after 74.07407407407408us,
    X"3df3b5" after 74.27427427427428us,
    X"3e76c8" after 74.47447447447448us,
    X"3ef9da" after 74.67467467467468us,
    X"3f7ced" after 74.87487487487488us,
    X"3fffff" after 75.07507507507508us,
    X"408311" after 75.27527527527528us,
    X"410624" after 75.47547547547548us,
    X"418936" after 75.67567567567568us,
    X"420c49" after 75.87587587587588us,
    X"428f5b" after 76.07607607607608us,
    X"43126e" after 76.27627627627628us,
    X"439580" after 76.47647647647648us,
    X"441892" after 76.67667667667668us,
    X"449ba5" after 76.87687687687688us,
    X"451eb7" after 77.07707707707708us,
    X"45a1ca" after 77.27727727727728us,
    X"4624dc" after 77.47747747747748us,
    X"46a7ef" after 77.67767767767768us,
    X"472b01" after 77.87787787787788us,
    X"47ae13" after 78.07807807807808us,
    X"483126" after 78.27827827827828us,
    X"48b438" after 78.47847847847848us,
    X"49374b" after 78.67867867867868us,
    X"49ba5d" after 78.87887887887888us,
    X"4a3d70" after 79.07907907907908us,
    X"4ac082" after 79.27927927927928us,
    X"4b4394" after 79.47947947947948us,
    X"4bc6a7" after 79.67967967967968us,
    X"4c49b9" after 79.87987987987988us,
    X"4ccccc" after 80.08008008008008us,
    X"4d4fde" after 80.28028028028028us,
    X"4dd2f1" after 80.48048048048048us,
    X"4e5603" after 80.68068068068068us,
    X"4ed915" after 80.88088088088088us,
    X"4f5c28" after 81.08108108108108us,
    X"4fdf3a" after 81.28128128128128us,
    X"50624d" after 81.48148148148148us,
    X"50e55f" after 81.68168168168168us,
    X"516872" after 81.88188188188188us,
    X"51eb84" after 82.08208208208208us,
    X"526e96" after 82.28228228228228us,
    X"52f1a9" after 82.48248248248248us,
    X"5374bb" after 82.68268268268268us,
    X"53f7ce" after 82.88288288288288us,
    X"547ae0" after 83.08308308308308us,
    X"54fdf3" after 83.28328328328328us,
    X"558105" after 83.48348348348348us,
    X"560417" after 83.68368368368368us,
    X"56872a" after 83.88388388388388us,
    X"570a3c" after 84.08408408408408us,
    X"578d4f" after 84.28428428428428us,
    X"581061" after 84.48448448448448us,
    X"589374" after 84.68468468468468us,
    X"591686" after 84.88488488488488us,
    X"599998" after 85.08508508508508us,
    X"5a1cab" after 85.28528528528528us,
    X"5a9fbd" after 85.4854854854855us,
    X"5b22d0" after 85.6856856856857us,
    X"5ba5e2" after 85.8858858858859us,
    X"5c28f5" after 86.0860860860861us,
    X"5cac07" after 86.2862862862863us,
    X"5d2f19" after 86.4864864864865us,
    X"5db22c" after 86.6866866866867us,
    X"5e353e" after 86.8868868868869us,
    X"5eb851" after 87.0870870870871us,
    X"5f3b63" after 87.2872872872873us,
    X"5fbe76" after 87.4874874874875us,
    X"604188" after 87.6876876876877us,
    X"60c49a" after 87.8878878878879us,
    X"6147ad" after 88.0880880880881us,
    X"61cabf" after 88.2882882882883us,
    X"624dd2" after 88.4884884884885us,
    X"62d0e4" after 88.6886886886887us,
    X"6353f7" after 88.8888888888889us,
    X"63d709" after 89.0890890890891us,
    X"645a1b" after 89.2892892892893us,
    X"64dd2e" after 89.4894894894895us,
    X"656040" after 89.6896896896897us,
    X"65e353" after 89.8898898898899us,
    X"666665" after 90.0900900900901us,
    X"66e978" after 90.2902902902903us,
    X"676c8a" after 90.4904904904905us,
    X"67ef9c" after 90.6906906906907us,
    X"6872af" after 90.8908908908909us,
    X"68f5c1" after 91.0910910910911us,
    X"6978d4" after 91.2912912912913us,
    X"69fbe6" after 91.4914914914915us,
    X"6a7ef9" after 91.6916916916917us,
    X"6b020b" after 91.8918918918919us,
    X"6b851d" after 92.0920920920921us,
    X"6c0830" after 92.2922922922923us,
    X"6c8b42" after 92.4924924924925us,
    X"6d0e55" after 92.6926926926927us,
    X"6d9167" after 92.8928928928929us,
    X"6e147a" after 93.0930930930931us,
    X"6e978c" after 93.2932932932933us,
    X"6f1a9e" after 93.4934934934935us,
    X"6f9db1" after 93.6936936936937us,
    X"7020c3" after 93.8938938938939us,
    X"70a3d6" after 94.0940940940941us,
    X"7126e8" after 94.2942942942943us,
    X"71a9fb" after 94.4944944944945us,
    X"722d0d" after 94.6946946946947us,
    X"72b01f" after 94.8948948948949us,
    X"733332" after 95.0950950950951us,
    X"73b644" after 95.2952952952953us,
    X"743957" after 95.4954954954955us,
    X"74bc69" after 95.6956956956957us,
    X"753f7c" after 95.8958958958959us,
    X"75c28e" after 96.0960960960961us,
    X"7645a0" after 96.2962962962963us,
    X"76c8b3" after 96.4964964964965us,
    X"774bc5" after 96.6966966966967us,
    X"77ced8" after 96.8968968968969us,
    X"7851ea" after 97.0970970970971us,
    X"78d4fd" after 97.2972972972973us,
    X"79580f" after 97.4974974974975us,
    X"79db21" after 97.6976976976977us,
    X"7a5e34" after 97.8978978978979us,
    X"7ae146" after 98.0980980980981us,
    X"7b6459" after 98.2982982982983us,
    X"7be76b" after 98.4984984984985us,
    X"7c6a7e" after 98.6986986986987us,
    X"7ced90" after 98.8988988988989us,
    X"7d70a2" after 99.0990990990991us,
    X"7df3b5" after 99.2992992992993us,
    X"7e76c7" after 99.4994994994995us,
    X"7ef9da" after 99.6996996996997us,
    X"7f7cec" after 99.8998998998999us,
    X"7fffff" after 100.10010010010011us,
    X"7f7cec" after 100.30030030030031us,
    X"7ef9da" after 100.50050050050051us,
    X"7e76c7" after 100.70070070070071us,
    X"7df3b5" after 100.90090090090091us,
    X"7d70a2" after 101.10110110110111us,
    X"7ced90" after 101.30130130130131us,
    X"7c6a7e" after 101.50150150150151us,
    X"7be76b" after 101.70170170170171us,
    X"7b6459" after 101.90190190190191us,
    X"7ae146" after 102.10210210210211us,
    X"7a5e34" after 102.30230230230231us,
    X"79db21" after 102.50250250250251us,
    X"79580f" after 102.70270270270271us,
    X"78d4fd" after 102.90290290290291us,
    X"7851ea" after 103.10310310310311us,
    X"77ced8" after 103.30330330330331us,
    X"774bc5" after 103.50350350350351us,
    X"76c8b3" after 103.70370370370371us,
    X"7645a0" after 103.90390390390391us,
    X"75c28e" after 104.10410410410411us,
    X"753f7c" after 104.30430430430431us,
    X"74bc69" after 104.50450450450451us,
    X"743957" after 104.70470470470471us,
    X"73b644" after 104.90490490490491us,
    X"733332" after 105.10510510510511us,
    X"72b01f" after 105.30530530530531us,
    X"722d0d" after 105.50550550550551us,
    X"71a9fb" after 105.70570570570571us,
    X"7126e8" after 105.90590590590591us,
    X"70a3d6" after 106.10610610610611us,
    X"7020c3" after 106.30630630630631us,
    X"6f9db1" after 106.50650650650651us,
    X"6f1a9e" after 106.70670670670671us,
    X"6e978c" after 106.90690690690691us,
    X"6e147a" after 107.10710710710711us,
    X"6d9167" after 107.30730730730731us,
    X"6d0e55" after 107.50750750750751us,
    X"6c8b42" after 107.70770770770771us,
    X"6c0830" after 107.90790790790791us,
    X"6b851d" after 108.10810810810811us,
    X"6b020b" after 108.30830830830831us,
    X"6a7ef9" after 108.50850850850851us,
    X"69fbe6" after 108.70870870870871us,
    X"6978d4" after 108.90890890890891us,
    X"68f5c1" after 109.10910910910911us,
    X"6872af" after 109.30930930930931us,
    X"67ef9c" after 109.50950950950951us,
    X"676c8a" after 109.70970970970971us,
    X"66e978" after 109.90990990990991us,
    X"666665" after 110.11011011011011us,
    X"65e353" after 110.31031031031031us,
    X"656040" after 110.51051051051051us,
    X"64dd2e" after 110.71071071071071us,
    X"645a1b" after 110.91091091091091us,
    X"63d709" after 111.11111111111111us,
    X"6353f7" after 111.31131131131131us,
    X"62d0e4" after 111.51151151151151us,
    X"624dd2" after 111.71171171171171us,
    X"61cabf" after 111.91191191191191us,
    X"6147ad" after 112.11211211211211us,
    X"60c49a" after 112.31231231231232us,
    X"604188" after 112.51251251251252us,
    X"5fbe76" after 112.71271271271272us,
    X"5f3b63" after 112.91291291291292us,
    X"5eb851" after 113.11311311311312us,
    X"5e353e" after 113.31331331331332us,
    X"5db22c" after 113.51351351351352us,
    X"5d2f19" after 113.71371371371372us,
    X"5cac07" after 113.91391391391392us,
    X"5c28f5" after 114.11411411411412us,
    X"5ba5e2" after 114.31431431431432us,
    X"5b22d0" after 114.51451451451452us,
    X"5a9fbd" after 114.71471471471472us,
    X"5a1cab" after 114.91491491491492us,
    X"599998" after 115.11511511511512us,
    X"591686" after 115.31531531531532us,
    X"589374" after 115.51551551551552us,
    X"581061" after 115.71571571571572us,
    X"578d4f" after 115.91591591591592us,
    X"570a3c" after 116.11611611611612us,
    X"56872a" after 116.31631631631632us,
    X"560417" after 116.51651651651652us,
    X"558105" after 116.71671671671672us,
    X"54fdf3" after 116.91691691691692us,
    X"547ae0" after 117.11711711711712us,
    X"53f7ce" after 117.31731731731732us,
    X"5374bb" after 117.51751751751752us,
    X"52f1a9" after 117.71771771771772us,
    X"526e96" after 117.91791791791792us,
    X"51eb84" after 118.11811811811812us,
    X"516872" after 118.31831831831832us,
    X"50e55f" after 118.51851851851852us,
    X"50624d" after 118.71871871871872us,
    X"4fdf3a" after 118.91891891891892us,
    X"4f5c28" after 119.11911911911912us,
    X"4ed915" after 119.31931931931932us,
    X"4e5603" after 119.51951951951952us,
    X"4dd2f1" after 119.71971971971973us,
    X"4d4fde" after 119.91991991991993us,
    X"4ccccc" after 120.12012012012013us,
    X"4c49b9" after 120.32032032032033us,
    X"4bc6a7" after 120.52052052052053us,
    X"4b4394" after 120.72072072072073us,
    X"4ac082" after 120.92092092092093us,
    X"4a3d70" after 121.12112112112113us,
    X"49ba5d" after 121.32132132132134us,
    X"49374b" after 121.52152152152154us,
    X"48b438" after 121.72172172172174us,
    X"483126" after 121.92192192192194us,
    X"47ae13" after 122.12212212212214us,
    X"472b01" after 122.32232232232234us,
    X"46a7ef" after 122.52252252252254us,
    X"4624dc" after 122.72272272272274us,
    X"45a1ca" after 122.92292292292294us,
    X"451eb7" after 123.12312312312314us,
    X"449ba5" after 123.32332332332334us,
    X"441892" after 123.52352352352354us,
    X"439580" after 123.72372372372374us,
    X"43126e" after 123.92392392392394us,
    X"428f5b" after 124.12412412412414us,
    X"420c49" after 124.32432432432434us,
    X"418936" after 124.52452452452454us,
    X"410624" after 124.72472472472474us,
    X"408311" after 124.92492492492494us,
    X"3fffff" after 125.12512512512514us,
    X"3f7ced" after 125.32532532532534us,
    X"3ef9da" after 125.52552552552554us,
    X"3e76c8" after 125.72572572572574us,
    X"3df3b5" after 125.92592592592594us,
    X"3d70a3" after 126.12612612612614us,
    X"3ced90" after 126.32632632632634us,
    X"3c6a7e" after 126.52652652652654us,
    X"3be76c" after 126.72672672672674us,
    X"3b6459" after 126.92692692692694us,
    X"3ae147" after 127.12712712712714us,
    X"3a5e34" after 127.32732732732734us,
    X"39db22" after 127.52752752752754us,
    X"39580f" after 127.72772772772774us,
    X"38d4fd" after 127.92792792792794us,
    X"3851eb" after 128.12812812812814us,
    X"37ced8" after 128.32832832832833us,
    X"374bc6" after 128.52852852852854us,
    X"36c8b3" after 128.72872872872873us,
    X"3645a1" after 128.92892892892894us,
    X"35c28e" after 129.12912912912913us,
    X"353f7c" after 129.32932932932934us,
    X"34bc6a" after 129.52952952952953us,
    X"343957" after 129.72972972972974us,
    X"33b645" after 129.92992992992993us,
    X"333332" after 130.13013013013014us,
    X"32b020" after 130.33033033033033us,
    X"322d0d" after 130.53053053053054us,
    X"31a9fb" after 130.73073073073073us,
    X"3126e9" after 130.93093093093094us,
    X"30a3d6" after 131.13113113113113us,
    X"3020c4" after 131.33133133133134us,
    X"2f9db1" after 131.53153153153153us,
    X"2f1a9f" after 131.73173173173174us,
    X"2e978c" after 131.93193193193193us,
    X"2e147a" after 132.13213213213214us,
    X"2d9168" after 132.33233233233233us,
    X"2d0e55" after 132.53253253253254us,
    X"2c8b43" after 132.73273273273273us,
    X"2c0830" after 132.93293293293294us,
    X"2b851e" after 133.13313313313313us,
    X"2b020b" after 133.33333333333334us,
    X"2a7ef9" after 133.53353353353353us,
    X"29fbe7" after 133.73373373373374us,
    X"2978d4" after 133.93393393393393us,
    X"28f5c2" after 134.13413413413414us,
    X"2872af" after 134.33433433433433us,
    X"27ef9d" after 134.53453453453454us,
    X"276c8a" after 134.73473473473473us,
    X"26e978" after 134.93493493493494us,
    X"266666" after 135.13513513513513us,
    X"25e353" after 135.33533533533534us,
    X"256041" after 135.53553553553553us,
    X"24dd2e" after 135.73573573573574us,
    X"245a1c" after 135.93593593593593us,
    X"23d709" after 136.13613613613614us,
    X"2353f7" after 136.33633633633633us,
    X"22d0e5" after 136.53653653653654us,
    X"224dd2" after 136.73673673673676us,
    X"21cac0" after 136.93693693693695us,
    X"2147ad" after 137.13713713713716us,
    X"20c49b" after 137.33733733733735us,
    X"204188" after 137.53753753753756us,
    X"1fbe76" after 137.73773773773775us,
    X"1f3b64" after 137.93793793793796us,
    X"1eb851" after 138.13813813813815us,
    X"1e353f" after 138.33833833833836us,
    X"1db22c" after 138.53853853853855us,
    X"1d2f1a" after 138.73873873873876us,
    X"1cac07" after 138.93893893893895us,
    X"1c28f5" after 139.13913913913916us,
    X"1ba5e3" after 139.33933933933935us,
    X"1b22d0" after 139.53953953953956us,
    X"1a9fbe" after 139.73973973973975us,
    X"1a1cab" after 139.93993993993996us,
    X"199999" after 140.14014014014015us,
    X"191686" after 140.34034034034036us,
    X"189374" after 140.54054054054055us,
    X"181062" after 140.74074074074076us,
    X"178d4f" after 140.94094094094095us,
    X"170a3d" after 141.14114114114116us,
    X"16872a" after 141.34134134134135us,
    X"160418" after 141.54154154154156us,
    X"158105" after 141.74174174174175us,
    X"14fdf3" after 141.94194194194196us,
    X"147ae1" after 142.14214214214215us,
    X"13f7ce" after 142.34234234234236us,
    X"1374bc" after 142.54254254254255us,
    X"12f1a9" after 142.74274274274276us,
    X"126e97" after 142.94294294294295us,
    X"11eb84" after 143.14314314314316us,
    X"116872" after 143.34334334334335us,
    X"10e560" after 143.54354354354356us,
    X"10624d" after 143.74374374374375us,
    X"0fdf3b" after 143.94394394394396us,
    X"0f5c28" after 144.14414414414415us,
    X"0ed916" after 144.34434434434436us,
    X"0e5603" after 144.54454454454455us,
    X"0dd2f1" after 144.74474474474476us,
    X"0d4fdf" after 144.94494494494495us,
    X"0ccccc" after 145.14514514514516us,
    X"0c49ba" after 145.34534534534535us,
    X"0bc6a7" after 145.54554554554556us,
    X"0b4395" after 145.74574574574575us,
    X"0ac082" after 145.94594594594597us,
    X"0a3d70" after 146.14614614614615us,
    X"09ba5e" after 146.34634634634637us,
    X"09374b" after 146.54654654654655us,
    X"08b439" after 146.74674674674677us,
    X"083126" after 146.94694694694695us,
    X"07ae14" after 147.14714714714717us,
    X"072b01" after 147.34734734734735us,
    X"06a7ef" after 147.54754754754757us,
    X"0624dd" after 147.74774774774775us,
    X"05a1ca" after 147.94794794794797us,
    X"051eb8" after 148.14814814814815us,
    X"049ba5" after 148.34834834834837us,
    X"041893" after 148.54854854854855us,
    X"039580" after 148.74874874874877us,
    X"03126e" after 148.94894894894895us,
    X"028f5c" after 149.14914914914917us,
    X"020c49" after 149.34934934934935us,
    X"018937" after 149.54954954954957us,
    X"010624" after 149.74974974974975us,
    X"008312" after 149.94994994994997us,
    X"ffffff" after 150.15015015015015us,
    X"ff7cec" after 150.35035035035037us,
    X"fef9da" after 150.55055055055055us,
    X"fe76c7" after 150.75075075075077us,
    X"fdf3b5" after 150.95095095095095us,
    X"fd70a2" after 151.15115115115117us,
    X"fced90" after 151.35135135135135us,
    X"fc6a7d" after 151.55155155155157us,
    X"fbe76b" after 151.75175175175175us,
    X"fb6459" after 151.95195195195197us,
    X"fae146" after 152.15215215215215us,
    X"fa5e34" after 152.35235235235237us,
    X"f9db21" after 152.55255255255256us,
    X"f9580f" after 152.75275275275277us,
    X"f8d4fc" after 152.95295295295296us,
    X"f851ea" after 153.15315315315317us,
    X"f7ced8" after 153.35335335335336us,
    X"f74bc5" after 153.55355355355357us,
    X"f6c8b3" after 153.75375375375376us,
    X"f645a0" after 153.95395395395397us,
    X"f5c28e" after 154.15415415415416us,
    X"f53f7b" after 154.35435435435437us,
    X"f4bc69" after 154.55455455455456us,
    X"f43957" after 154.75475475475477us,
    X"f3b644" after 154.95495495495496us,
    X"f33332" after 155.15515515515517us,
    X"f2b01f" after 155.35535535535536us,
    X"f22d0d" after 155.55555555555557us,
    X"f1a9fa" after 155.75575575575576us,
    X"f126e8" after 155.95595595595597us,
    X"f0a3d6" after 156.15615615615616us,
    X"f020c3" after 156.35635635635637us,
    X"ef9db1" after 156.55655655655656us,
    X"ef1a9e" after 156.75675675675677us,
    X"ee978c" after 156.95695695695696us,
    X"ee1479" after 157.15715715715717us,
    X"ed9167" after 157.35735735735736us,
    X"ed0e55" after 157.55755755755757us,
    X"ec8b42" after 157.75775775775776us,
    X"ec0830" after 157.95795795795797us,
    X"eb851d" after 158.15815815815816us,
    X"eb020b" after 158.35835835835837us,
    X"ea7ef8" after 158.55855855855856us,
    X"e9fbe6" after 158.75875875875877us,
    X"e978d3" after 158.95895895895896us,
    X"e8f5c1" after 159.15915915915917us,
    X"e872af" after 159.35935935935936us,
    X"e7ef9c" after 159.55955955955957us,
    X"e76c8a" after 159.75975975975976us,
    X"e6e977" after 159.95995995995997us,
    X"e66665" after 160.16016016016016us,
    X"e5e352" after 160.36036036036037us,
    X"e56040" after 160.56056056056056us,
    X"e4dd2e" after 160.76076076076077us,
    X"e45a1b" after 160.96096096096096us,
    X"e3d709" after 161.16116116116117us,
    X"e353f6" after 161.36136136136136us,
    X"e2d0e4" after 161.56156156156158us,
    X"e24dd1" after 161.76176176176176us,
    X"e1cabf" after 161.96196196196198us,
    X"e147ad" after 162.16216216216216us,
    X"e0c49a" after 162.36236236236238us,
    X"e04188" after 162.56256256256256us,
    X"dfbe75" after 162.76276276276278us,
    X"df3b63" after 162.96296296296296us,
    X"deb850" after 163.16316316316318us,
    X"de353e" after 163.36336336336336us,
    X"ddb22c" after 163.56356356356358us,
    X"dd2f19" after 163.76376376376376us,
    X"dcac07" after 163.96396396396398us,
    X"dc28f4" after 164.16416416416416us,
    X"dba5e2" after 164.36436436436438us,
    X"db22cf" after 164.56456456456456us,
    X"da9fbd" after 164.76476476476478us,
    X"da1cab" after 164.96496496496496us,
    X"d99998" after 165.16516516516518us,
    X"d91686" after 165.36536536536536us,
    X"d89373" after 165.56556556556558us,
    X"d81061" after 165.76576576576576us,
    X"d78d4e" after 165.96596596596598us,
    X"d70a3c" after 166.16616616616616us,
    X"d6872a" after 166.36636636636638us,
    X"d60417" after 166.56656656656656us,
    X"d58105" after 166.76676676676678us,
    X"d4fdf2" after 166.96696696696696us,
    X"d47ae0" after 167.16716716716718us,
    X"d3f7cd" after 167.36736736736736us,
    X"d374bb" after 167.56756756756758us,
    X"d2f1a8" after 167.76776776776777us,
    X"d26e96" after 167.96796796796798us,
    X"d1eb84" after 168.16816816816817us,
    X"d16871" after 168.36836836836838us,
    X"d0e55f" after 168.56856856856857us,
    X"d0624c" after 168.76876876876878us,
    X"cfdf3a" after 168.96896896896897us,
    X"cf5c27" after 169.16916916916918us,
    X"ced915" after 169.36936936936937us,
    X"ce5603" after 169.56956956956958us,
    X"cdd2f0" after 169.76976976976977us,
    X"cd4fde" after 169.96996996996998us,
    X"cccccb" after 170.17017017017017us,
    X"cc49b9" after 170.37037037037038us,
    X"cbc6a6" after 170.57057057057057us,
    X"cb4394" after 170.77077077077078us,
    X"cac082" after 170.970970970971us,
    X"ca3d6f" after 171.17117117117118us,
    X"c9ba5d" after 171.3713713713714us,
    X"c9374a" after 171.57157157157158us,
    X"c8b438" after 171.7717717717718us,
    X"c83125" after 171.97197197197198us,
    X"c7ae13" after 172.1721721721722us,
    X"c72b01" after 172.37237237237238us,
    X"c6a7ee" after 172.5725725725726us,
    X"c624dc" after 172.77277277277278us,
    X"c5a1c9" after 172.972972972973us,
    X"c51eb7" after 173.17317317317318us,
    X"c49ba4" after 173.3733733733734us,
    X"c41892" after 173.57357357357358us,
    X"c39580" after 173.7737737737738us,
    X"c3126d" after 173.97397397397398us,
    X"c28f5b" after 174.1741741741742us,
    X"c20c48" after 174.37437437437438us,
    X"c18936" after 174.5745745745746us,
    X"c10623" after 174.77477477477478us,
    X"c08311" after 174.974974974975us,
    X"bfffff" after 175.17517517517518us,
    X"bf7cec" after 175.3753753753754us,
    X"bef9da" after 175.57557557557558us,
    X"be76c7" after 175.7757757757758us,
    X"bdf3b5" after 175.97597597597598us,
    X"bd70a2" after 176.1761761761762us,
    X"bced90" after 176.37637637637638us,
    X"bc6a7d" after 176.5765765765766us,
    X"bbe76b" after 176.77677677677679us,
    X"bb6459" after 176.976976976977us,
    X"bae146" after 177.17717717717719us,
    X"ba5e34" after 177.3773773773774us,
    X"b9db21" after 177.57757757757759us,
    X"b9580f" after 177.7777777777778us,
    X"b8d4fc" after 177.977977977978us,
    X"b851ea" after 178.1781781781782us,
    X"b7ced8" after 178.3783783783784us,
    X"b74bc5" after 178.5785785785786us,
    X"b6c8b3" after 178.7787787787788us,
    X"b645a0" after 178.978978978979us,
    X"b5c28e" after 179.1791791791792us,
    X"b53f7b" after 179.3793793793794us,
    X"b4bc69" after 179.5795795795796us,
    X"b43957" after 179.7797797797798us,
    X"b3b644" after 179.97997997998us,
    X"b33332" after 180.1801801801802us,
    X"b2b01f" after 180.3803803803804us,
    X"b22d0d" after 180.5805805805806us,
    X"b1a9fa" after 180.7807807807808us,
    X"b126e8" after 180.980980980981us,
    X"b0a3d6" after 181.1811811811812us,
    X"b020c3" after 181.3813813813814us,
    X"af9db1" after 181.5815815815816us,
    X"af1a9e" after 181.7817817817818us,
    X"ae978c" after 181.981981981982us,
    X"ae1479" after 182.1821821821822us,
    X"ad9167" after 182.3823823823824us,
    X"ad0e55" after 182.5825825825826us,
    X"ac8b42" after 182.7827827827828us,
    X"ac0830" after 182.982982982983us,
    X"ab851d" after 183.1831831831832us,
    X"ab020b" after 183.3833833833834us,
    X"aa7ef8" after 183.5835835835836us,
    X"a9fbe6" after 183.7837837837838us,
    X"a978d3" after 183.983983983984us,
    X"a8f5c1" after 184.1841841841842us,
    X"a872af" after 184.3843843843844us,
    X"a7ef9c" after 184.5845845845846us,
    X"a76c8a" after 184.7847847847848us,
    X"a6e977" after 184.984984984985us,
    X"a66665" after 185.1851851851852us,
    X"a5e352" after 185.3853853853854us,
    X"a56040" after 185.5855855855856us,
    X"a4dd2e" after 185.7857857857858us,
    X"a45a1b" after 185.985985985986us,
    X"a3d709" after 186.1861861861862us,
    X"a353f6" after 186.3863863863864us,
    X"a2d0e4" after 186.5865865865866us,
    X"a24dd1" after 186.7867867867868us,
    X"a1cabf" after 186.986986986987us,
    X"a147ad" after 187.1871871871872us,
    X"a0c49a" after 187.3873873873874us,
    X"a04188" after 187.5875875875876us,
    X"9fbe75" after 187.7877877877878us,
    X"9f3b63" after 187.987987987988us,
    X"9eb850" after 188.1881881881882us,
    X"9e353e" after 188.3883883883884us,
    X"9db22c" after 188.5885885885886us,
    X"9d2f19" after 188.7887887887888us,
    X"9cac07" after 188.988988988989us,
    X"9c28f4" after 189.1891891891892us,
    X"9ba5e2" after 189.3893893893894us,
    X"9b22cf" after 189.5895895895896us,
    X"9a9fbd" after 189.7897897897898us,
    X"9a1cab" after 189.98998998999us,
    X"999998" after 190.1901901901902us,
    X"991686" after 190.3903903903904us,
    X"989373" after 190.5905905905906us,
    X"981061" after 190.7907907907908us,
    X"978d4e" after 190.990990990991us,
    X"970a3c" after 191.1911911911912us,
    X"96872a" after 191.3913913913914us,
    X"960417" after 191.5915915915916us,
    X"958105" after 191.7917917917918us,
    X"94fdf2" after 191.991991991992us,
    X"947ae0" after 192.1921921921922us,
    X"93f7cd" after 192.3923923923924us,
    X"9374bb" after 192.5925925925926us,
    X"92f1a8" after 192.7927927927928us,
    X"926e96" after 192.992992992993us,
    X"91eb84" after 193.1931931931932us,
    X"916871" after 193.3933933933934us,
    X"90e55f" after 193.5935935935936us,
    X"90624c" after 193.7937937937938us,
    X"8fdf3a" after 193.993993993994us,
    X"8f5c27" after 194.1941941941942us,
    X"8ed915" after 194.3943943943944us,
    X"8e5603" after 194.5945945945946us,
    X"8dd2f0" after 194.7947947947948us,
    X"8d4fde" after 194.994994994995us,
    X"8ccccb" after 195.1951951951952us,
    X"8c49b9" after 195.3953953953954us,
    X"8bc6a6" after 195.5955955955956us,
    X"8b4394" after 195.7957957957958us,
    X"8ac082" after 195.995995995996us,
    X"8a3d6f" after 196.1961961961962us,
    X"89ba5d" after 196.3963963963964us,
    X"89374a" after 196.5965965965966us,
    X"88b438" after 196.7967967967968us,
    X"883125" after 196.996996996997us,
    X"87ae13" after 197.1971971971972us,
    X"872b01" after 197.3973973973974us,
    X"86a7ee" after 197.5975975975976us,
    X"8624dc" after 197.7977977977978us,
    X"85a1c9" after 197.997997997998us,
    X"851eb7" after 198.1981981981982us,
    X"849ba4" after 198.3983983983984us,
    X"841892" after 198.5985985985986us,
    X"839580" after 198.7987987987988us,
    X"83126d" after 198.998998998999us,
    X"828f5b" after 199.1991991991992us,
    X"820c48" after 199.3993993993994us,
    X"818936" after 199.5995995995996us,
    X"810623" after 199.7997997997998us,
    X"808311" after 200.0us;
    
    -- etude en NAND
    /*Vin <= X"ffffffff" after 0.0us,
    X"ffffffff" after 0.10005002501250625us,
    X"ffffffff" after 0.2001000500250125us,
    X"ffffffff" after 0.3001500750375187us,
    X"ffffffff" after 0.400200100050025us,
    X"ffffffff" after 0.5002501250625312us,
    X"ffffffff" after 0.6003001500750375us,
    X"ffffffff" after 0.7003501750875437us,
    X"ffffffff" after 0.80040020010005us,
    X"ffffffff" after 0.9004502251125562us,
    X"ffffffff" after 1.0005002501250624us,
    X"ffffffff" after 1.1005502751375686us,
    X"ffffffff" after 1.200600300150075us,
    X"ffffffff" after 1.3006503251625812us,
    X"ffffffff" after 1.4007003501750874us,
    X"ffffffff" after 1.5007503751875937us,
    X"ffffffff" after 1.6008004002001us,
    X"ffffffff" after 1.7008504252126062us,
    X"ffffffff" after 1.8009004502251125us,
    X"ffffffff" after 1.9009504752376187us,
    X"ffffffff" after 2.0010005002501248us,
    X"ffffffff" after 2.101050525262631us,
    X"ffffffff" after 2.2011005502751373us,
    X"ffffffff" after 2.3011505752876436us,
    X"ffffffff" after 2.40120060030015us,
    X"ffffffff" after 2.501250625312656us,
    X"ffffffff" after 2.6013006503251623us,
    X"ffffffff" after 2.7013506753376686us,
    X"ffffffff" after 2.801400700350175us,
    X"ffffffff" after 2.901450725362681us,
    X"ffffffff" after 3.0015007503751874us,
    X"ffffffff" after 3.1015507753876936us,
    X"ffffffff" after 3.2016008004002us,
    X"ffffffff" after 3.301650825412706us,
    X"ffffffff" after 3.4017008504252124us,
    X"ffffffff" after 3.5017508754377187us,
    X"ffffffff" after 3.601800900450225us,
    X"ffffffff" after 3.701850925462731us,
    X"ffffffff" after 3.8019009504752375us,
    X"ffffffff" after 3.9019509754877437us,
    X"ffffffff" after 4.0020010005002495us,
    X"ffffffff" after 4.102051025512756us,
    X"ffffffff" after 4.202101050525262us,
    X"ffffffff" after 4.302151075537768us,
    X"ffffffff" after 4.402201100550275us,
    X"ffffffff" after 4.502251125562781us,
    X"ffffffff" after 4.602301150575287us,
    X"ffffffff" after 4.702351175587793us,
    X"ffffffff" after 4.8024012006003us,
    X"ffffffff" after 4.902451225612806us,
    X"80000000" after 5.002501250625312us,
    X"80000000" after 5.102551275637818us,
    X"80000000" after 5.202601300650325us,
    X"80000000" after 5.302651325662831us,
    X"80000000" after 5.402701350675337us,
    X"80000000" after 5.5027513756878434us,
    X"80000000" after 5.60280140070035us,
    X"80000000" after 5.702851425712856us,
    X"80000000" after 5.802901450725362us,
    X"80000000" after 5.9029514757378685us,
    X"80000000" after 6.003001500750375us,
    X"80000000" after 6.103051525762881us,
    X"80000000" after 6.203101550775387us,
    X"80000000" after 6.3031515757878935us,
    X"80000000" after 6.4032016008004us,
    X"80000000" after 6.503251625812906us,
    X"80000000" after 6.603301650825412us,
    X"80000000" after 6.703351675837919us,
    X"80000000" after 6.803401700850425us,
    X"80000000" after 6.903451725862931us,
    X"80000000" after 7.003501750875437us,
    X"80000000" after 7.103551775887944us,
    X"80000000" after 7.20360180090045us,
    X"80000000" after 7.303651825912956us,
    X"80000000" after 7.403701850925462us,
    X"80000000" after 7.503751875937969us,
    X"80000000" after 7.603801900950475us,
    X"80000000" after 7.703851925962981us,
    X"80000000" after 7.8039019509754874us,
    X"80000000" after 7.903951975987994us,
    X"80000000" after 8.004002001000499us,
    X"80000000" after 8.104052026013006us,
    X"80000000" after 8.204102051025512us,
    X"80000000" after 8.304152076038019us,
    X"80000000" after 8.404202101050524us,
    X"80000000" after 8.504252126063031us,
    X"80000000" after 8.604302151075537us,
    X"80000000" after 8.704352176088044us,
    X"80000000" after 8.80440220110055us,
    X"80000000" after 8.904452226113056us,
    X"80000000" after 9.004502251125562us,
    X"80000000" after 9.104552276138069us,
    X"80000000" after 9.204602301150574us,
    X"80000000" after 9.304652326163081us,
    X"80000000" after 9.404702351175587us,
    X"80000000" after 9.504752376188094us,
    X"80000000" after 9.6048024012006us,
    X"80000000" after 9.704852426213106us,
    X"80000000" after 9.804902451225612us,
    X"80000000" after 9.904952476238119us,
    X"80000000" after 10.005002501250624us,
    X"80000000" after 10.105052526263131us,
    X"80000000" after 10.205102551275637us,
    X"80000000" after 10.305152576288144us,
    X"80000000" after 10.40520260130065us,
    X"80000000" after 10.505252626313156us,
    X"80000000" after 10.605302651325662us,
    X"80000000" after 10.705352676338169us,
    X"80000000" after 10.805402701350674us,
    X"80000000" after 10.905452726363182us,
    X"80000000" after 11.005502751375687us,
    X"80000000" after 11.105552776388194us,
    X"80000000" after 11.2056028014007us,
    X"80000000" after 11.305652826413207us,
    X"80000000" after 11.405702851425712us,
    X"80000000" after 11.505752876438219us,
    X"80000000" after 11.605802901450724us,
    X"80000000" after 11.705852926463232us,
    X"80000000" after 11.805902951475737us,
    X"80000000" after 11.905952976488244us,
    X"80000000" after 12.00600300150075us,
    X"80000000" after 12.106053026513257us,
    X"80000000" after 12.206103051525762us,
    X"80000000" after 12.30615307653827us,
    X"80000000" after 12.406203101550775us,
    X"80000000" after 12.506253126563282us,
    X"80000000" after 12.606303151575787us,
    X"80000000" after 12.706353176588294us,
    X"80000000" after 12.8064032016008us,
    X"80000000" after 12.906453226613305us,
    X"80000000" after 13.006503251625812us,
    X"80000000" after 13.106553276638317us,
    X"80000000" after 13.206603301650825us,
    X"80000000" after 13.30665332666333us,
    X"80000000" after 13.406703351675837us,
    X"80000000" after 13.506753376688343us,
    X"80000000" after 13.60680340170085us,
    X"80000000" after 13.706853426713355us,
    X"80000000" after 13.806903451725862us,
    X"80000000" after 13.906953476738368us,
    X"80000000" after 14.007003501750875us,
    X"80000000" after 14.10705352676338us,
    X"80000000" after 14.207103551775887us,
    X"80000000" after 14.307153576788393us,
    X"80000000" after 14.4072036018009us,
    X"80000000" after 14.507253626813405us,
    X"80000000" after 14.607303651825912us,
    X"80000000" after 14.707353676838418us,
    X"80000000" after 14.807403701850925us,
    X"80000000" after 14.90745372686343us,
    X"ffffffff" after 15.007503751875937us,
    X"ffffffff" after 15.107553776888443us,
    X"ffffffff" after 15.20760380190095us,
    X"ffffffff" after 15.307653826913455us,
    X"ffffffff" after 15.407703851925962us,
    X"ffffffff" after 15.507753876938468us,
    X"ffffffff" after 15.607803901950975us,
    X"ffffffff" after 15.70785392696348us,
    X"ffffffff" after 15.807903951975987us,
    X"ffffffff" after 15.907953976988493us,
    X"ffffffff" after 16.008004002000998us,
    X"ffffffff" after 16.108054027013505us,
    X"ffffffff" after 16.208104052026012us,
    X"ffffffff" after 16.30815407703852us,
    X"ffffffff" after 16.408204102051023us,
    X"ffffffff" after 16.50825412706353us,
    X"ffffffff" after 16.608304152076037us,
    X"ffffffff" after 16.708354177088545us,
    X"ffffffff" after 16.80840420210105us,
    X"ffffffff" after 16.908454227113555us,
    X"ffffffff" after 17.008504252126063us,
    X"ffffffff" after 17.10855427713857us,
    X"ffffffff" after 17.208604302151073us,
    X"ffffffff" after 17.30865432716358us,
    X"ffffffff" after 17.408704352176088us,
    X"ffffffff" after 17.508754377188595us,
    X"ffffffff" after 17.6088044022011us,
    X"ffffffff" after 17.708854427213605us,
    X"ffffffff" after 17.808904452226113us,
    X"ffffffff" after 17.90895447723862us,
    X"ffffffff" after 18.009004502251123us,
    X"ffffffff" after 18.10905452726363us,
    X"ffffffff" after 18.209104552276138us,
    X"ffffffff" after 18.309154577288645us,
    X"ffffffff" after 18.40920460230115us,
    X"ffffffff" after 18.509254627313656us,
    X"ffffffff" after 18.609304652326163us,
    X"ffffffff" after 18.70935467733867us,
    X"ffffffff" after 18.809404702351173us,
    X"ffffffff" after 18.90945472736368us,
    X"ffffffff" after 19.009504752376188us,
    X"ffffffff" after 19.109554777388695us,
    X"ffffffff" after 19.2096048024012us,
    X"ffffffff" after 19.309654827413706us,
    X"ffffffff" after 19.409704852426213us,
    X"ffffffff" after 19.509754877438716us,
    X"ffffffff" after 19.609804902451224us,
    X"ffffffff" after 19.70985492746373us,
    X"ffffffff" after 19.809904952476238us,
    X"ffffffff" after 19.90995497748874us,
    X"ffffffff" after 20.01000500250125us,
    X"ffffffff" after 20.110055027513756us,
    X"ffffffff" after 20.210105052526263us,
    X"ffffffff" after 20.310155077538766us,
    X"ffffffff" after 20.410205102551274us,
    X"ffffffff" after 20.51025512756378us,
    X"ffffffff" after 20.610305152576288us,
    X"ffffffff" after 20.71035517758879us,
    X"ffffffff" after 20.8104052026013us,
    X"ffffffff" after 20.910455227613806us,
    X"ffffffff" after 21.010505252626313us,
    X"ffffffff" after 21.110555277638817us,
    X"ffffffff" after 21.210605302651324us,
    X"ffffffff" after 21.31065532766383us,
    X"ffffffff" after 21.410705352676338us,
    X"ffffffff" after 21.51075537768884us,
    X"ffffffff" after 21.61080540270135us,
    X"ffffffff" after 21.710855427713856us,
    X"ffffffff" after 21.810905452726363us,
    X"ffffffff" after 21.910955477738867us,
    X"ffffffff" after 22.011005502751374us,
    X"ffffffff" after 22.11105552776388us,
    X"ffffffff" after 22.211105552776388us,
    X"ffffffff" after 22.31115557778889us,
    X"ffffffff" after 22.4112056028014us,
    X"ffffffff" after 22.511255627813906us,
    X"ffffffff" after 22.611305652826413us,
    X"ffffffff" after 22.711355677838917us,
    X"ffffffff" after 22.811405702851424us,
    X"ffffffff" after 22.91145572786393us,
    X"ffffffff" after 23.011505752876438us,
    X"ffffffff" after 23.11155577788894us,
    X"ffffffff" after 23.21160580290145us,
    X"ffffffff" after 23.311655827913956us,
    X"ffffffff" after 23.411705852926463us,
    X"ffffffff" after 23.511755877938967us,
    X"ffffffff" after 23.611805902951474us,
    X"ffffffff" after 23.71185592796398us,
    X"ffffffff" after 23.81190595297649us,
    X"ffffffff" after 23.911955977988992us,
    X"ffffffff" after 24.0120060030015us,
    X"ffffffff" after 24.112056028014006us,
    X"ffffffff" after 24.212106053026513us,
    X"ffffffff" after 24.312156078039017us,
    X"ffffffff" after 24.412206103051524us,
    X"ffffffff" after 24.51225612806403us,
    X"ffffffff" after 24.61230615307654us,
    X"ffffffff" after 24.712356178089042us,
    X"ffffffff" after 24.81240620310155us,
    X"ffffffff" after 24.912456228114056us,
    X"ffffffff" after 25.012506253126563us,
    X"ffffffff" after 25.112556278139067us,
    X"ffffffff" after 25.212606303151574us,
    X"ffffffff" after 25.31265632816408us,
    X"ffffffff" after 25.41270635317659us,
    X"ffffffff" after 25.512756378189092us,
    X"ffffffff" after 25.6128064032016us,
    X"ffffffff" after 25.712856428214106us,
    X"ffffffff" after 25.81290645322661us,
    X"ffffffff" after 25.912956478239117us,
    X"ffffffff" after 26.013006503251624us,
    X"ffffffff" after 26.11305652826413us,
    X"ffffffff" after 26.213106553276635us,
    X"ffffffff" after 26.313156578289142us,
    X"ffffffff" after 26.41320660330165us,
    X"ffffffff" after 26.513256628314156us,
    X"ffffffff" after 26.61330665332666us,
    X"ffffffff" after 26.713356678339167us,
    X"ffffffff" after 26.813406703351674us,
    X"ffffffff" after 26.91345672836418us,
    X"ffffffff" after 27.013506753376685us,
    X"ffffffff" after 27.113556778389192us,
    X"ffffffff" after 27.2136068034017us,
    X"ffffffff" after 27.313656828414207us,
    X"ffffffff" after 27.41370685342671us,
    X"ffffffff" after 27.513756878439217us,
    X"ffffffff" after 27.613806903451724us,
    X"ffffffff" after 27.71385692846423us,
    X"ffffffff" after 27.813906953476735us,
    X"ffffffff" after 27.913956978489242us,
    X"ffffffff" after 28.01400700350175us,
    X"ffffffff" after 28.114057028514257us,
    X"ffffffff" after 28.21410705352676us,
    X"ffffffff" after 28.314157078539267us,
    X"ffffffff" after 28.414207103551774us,
    X"ffffffff" after 28.51425712856428us,
    X"ffffffff" after 28.614307153576785us,
    X"ffffffff" after 28.714357178589292us,
    X"ffffffff" after 28.8144072036018us,
    X"ffffffff" after 28.914457228614307us,
    X"ffffffff" after 29.01450725362681us,
    X"ffffffff" after 29.114557278639317us,
    X"ffffffff" after 29.214607303651825us,
    X"ffffffff" after 29.31465732866433us,
    X"ffffffff" after 29.414707353676835us,
    X"ffffffff" after 29.514757378689342us,
    X"ffffffff" after 29.61480740370185us,
    X"ffffffff" after 29.714857428714357us,
    X"ffffffff" after 29.81490745372686us,
    X"ffffffff" after 29.914957478739368us,
    X"7f800000" after 30.015007503751875us,
    X"7f800000" after 30.115057528764382us,
    X"7f800000" after 30.215107553776885us,
    X"7f800000" after 30.315157578789393us,
    X"7f800000" after 30.4152076038019us,
    X"7f800000" after 30.515257628814407us,
    X"7f800000" after 30.61530765382691us,
    X"7f800000" after 30.715357678839418us,
    X"7f800000" after 30.815407703851925us,
    X"7f800000" after 30.915457728864432us,
    X"7f800000" after 31.015507753876935us,
    X"7f800000" after 31.115557778889443us,
    X"7f800000" after 31.21560780390195us,
    X"7f800000" after 31.315657828914457us,
    X"7f800000" after 31.41570785392696us,
    X"7f800000" after 31.515757878939468us,
    X"7f800000" after 31.615807903951975us,
    X"7f800000" after 31.715857928964482us,
    X"7f800000" after 31.815907953976986us,
    X"7f800000" after 31.915957978989493us,
    X"7f800000" after 32.016008004001996us,
    X"7f800000" after 32.1160580290145us,
    X"7f800000" after 32.21610805402701us,
    X"7f800000" after 32.31615807903952us,
    X"7f800000" after 32.416208104052025us,
    X"7f800000" after 32.51625812906453us,
    X"7f800000" after 32.61630815407704us,
    X"7f800000" after 32.71635817908954us,
    X"7f800000" after 32.816408204102046us,
    X"7f800000" after 32.91645822911455us,
    X"7f800000" after 33.01650825412706us,
    X"7f800000" after 33.11655827913957us,
    X"7f800000" after 33.216608304152075us,
    X"7f800000" after 33.31665832916458us,
    X"7f800000" after 33.41670835417709us,
    X"7f800000" after 33.51675837918959us,
    X"7f800000" after 33.6168084042021us,
    X"7f800000" after 33.716858429214604us,
    X"7f800000" after 33.81690845422711us,
    X"7f800000" after 33.91695847923962us,
    X"7f800000" after 34.017008504252125us,
    X"7f800000" after 34.11705852926463us,
    X"7f800000" after 34.21710855427714us,
    X"7f800000" after 34.31715857928964us,
    X"7f800000" after 34.41720860430215us,
    X"7f800000" after 34.517258629314654us,
    X"7f800000" after 34.61730865432716us,
    X"7f800000" after 34.71735867933967us,
    X"7f800000" after 34.817408704352175us,
    X"7f800000" after 34.91745872936468us,
    X"7f800000" after 35.01750875437719us,
    X"7f800000" after 35.11755877938969us,
    X"7f800000" after 35.2176088044022us,
    X"7f800000" after 35.317658829414704us,
    X"7f800000" after 35.41770885442721us,
    X"7f800000" after 35.51775887943972us,
    X"7f800000" after 35.617808904452225us,
    X"7f800000" after 35.71785892946473us,
    X"7f800000" after 35.81790895447724us,
    X"7f800000" after 35.91795897948974us,
    X"7f800000" after 36.01800900450225us,
    X"7f800000" after 36.118059029514754us,
    X"7f800000" after 36.21810905452726us,
    X"7f800000" after 36.31815907953977us,
    X"7f800000" after 36.418209104552275us,
    X"7f800000" after 36.51825912956478us,
    X"7f800000" after 36.61830915457729us,
    X"7f800000" after 36.71835917958979us,
    X"7f800000" after 36.8184092046023us,
    X"7f800000" after 36.918459229614804us,
    X"7f800000" after 37.01850925462731us,
    X"7f800000" after 37.11855927963982us,
    X"7f800000" after 37.218609304652325us,
    X"7f800000" after 37.31865932966483us,
    X"7f800000" after 37.41870935467734us,
    X"7f800000" after 37.51875937968984us,
    X"7f800000" after 37.61880940470235us,
    X"7f800000" after 37.718859429714854us,
    X"7f800000" after 37.81890945472736us,
    X"7f800000" after 37.91895947973987us,
    X"7f800000" after 38.019009504752376us,
    X"7f800000" after 38.11905952976488us,
    X"7f800000" after 38.21910955477739us,
    X"7f800000" after 38.31915957978989us,
    X"7f800000" after 38.4192096048024us,
    X"7f800000" after 38.519259629814904us,
    X"7f800000" after 38.61930965482741us,
    X"7f800000" after 38.71935967983992us,
    X"7f800000" after 38.819409704852426us,
    X"7f800000" after 38.91945972986493us,
    X"7f800000" after 39.01950975487743us,
    X"7f800000" after 39.11955977988994us,
    X"7f800000" after 39.21960980490245us,
    X"7f800000" after 39.319659829914954us,
    X"7f800000" after 39.41970985492746us,
    X"7f800000" after 39.51975987993997us,
    X"7f800000" after 39.619809904952476us,
    X"7f800000" after 39.71985992996498us,
    X"7f800000" after 39.81990995497748us,
    X"7f800000" after 39.91995997998999us,
    X"ffffffff" after 40.0200100050025us,
    X"ffffffff" after 40.120060030015004us,
    X"ffffffff" after 40.22011005502751us,
    X"ffffffff" after 40.32016008004002us,
    X"ffffffff" after 40.420210105052526us,
    X"ffffffff" after 40.52026013006503us,
    X"ffffffff" after 40.62031015507753us,
    X"ffffffff" after 40.72036018009004us,
    X"ffffffff" after 40.82041020510255us,
    X"ffffffff" after 40.920460230115054us,
    X"ffffffff" after 41.02051025512756us,
    X"ffffffff" after 41.12056028014007us,
    X"ffffffff" after 41.220610305152576us,
    X"ffffffff" after 41.32066033016508us,
    X"ffffffff" after 41.42071035517758us,
    X"ffffffff" after 41.52076038019009us,
    X"ffffffff" after 41.6208104052026us,
    X"ffffffff" after 41.720860430215104us,
    X"ffffffff" after 41.82091045522761us,
    X"ffffffff" after 41.92096048024012us,
    X"ffffffff" after 42.021010505252626us,
    X"ffffffff" after 42.12106053026513us,
    X"ffffffff" after 42.22111055527763us,
    X"ffffffff" after 42.32116058029014us,
    X"ffffffff" after 42.42121060530265us,
    X"ffffffff" after 42.521260630315155us,
    X"ffffffff" after 42.62131065532766us,
    X"ffffffff" after 42.72136068034017us,
    X"ffffffff" after 42.821410705352676us,
    X"ffffffff" after 42.92146073036518us,
    X"ffffffff" after 43.02151075537768us,
    X"ffffffff" after 43.12156078039019us,
    X"ffffffff" after 43.2216108054027us,
    X"ffffffff" after 43.321660830415205us,
    X"ffffffff" after 43.42171085542771us,
    X"ffffffff" after 43.52176088044022us,
    X"ffffffff" after 43.621810905452726us,
    X"ffffffff" after 43.72186093046523us,
    X"ffffffff" after 43.82191095547773us,
    X"ffffffff" after 43.92196098049024us,
    X"ffffffff" after 44.02201100550275us,
    X"ffffffff" after 44.122061030515255us,
    X"ffffffff" after 44.22211105552776us,
    X"ffffffff" after 44.32216108054027us,
    X"ffffffff" after 44.422211105552776us,
    X"ffffffff" after 44.52226113056528us,
    X"ffffffff" after 44.62231115557778us,
    X"ffffffff" after 44.72236118059029us,
    X"ffffffff" after 44.8224112056028us,
    X"ffffffff" after 44.922461230615305us,
    X"ffffffff" after 45.02251125562781us,
    X"ffffffff" after 45.12256128064032us,
    X"ffffffff" after 45.222611305652826us,
    X"ffffffff" after 45.322661330665326us,
    X"ffffffff" after 45.42271135567783us,
    X"ffffffff" after 45.52276138069034us,
    X"ffffffff" after 45.62281140570285us,
    X"ffffffff" after 45.722861430715355us,
    X"ffffffff" after 45.82291145572786us,
    X"ffffffff" after 45.92296148074037us,
    X"ffffffff" after 46.023011505752876us,
    X"ffffffff" after 46.123061530765376us,
    X"ffffffff" after 46.22311155577788us,
    X"ffffffff" after 46.32316158079039us,
    X"ffffffff" after 46.4232116058029us,
    X"ffffffff" after 46.523261630815405us,
    X"ffffffff" after 46.62331165582791us,
    X"ffffffff" after 46.72336168084042us,
    X"ffffffff" after 46.823411705852926us,
    X"ffffffff" after 46.92346173086543us,
    X"ffffffff" after 47.023511755877934us,
    X"ffffffff" after 47.12356178089044us,
    X"ffffffff" after 47.22361180590295us,
    X"ffffffff" after 47.323661830915455us,
    X"ffffffff" after 47.42371185592796us,
    X"ffffffff" after 47.52376188094047us,
    X"ffffffff" after 47.62381190595298us,
    X"ffffffff" after 47.72386193096548us,
    X"ffffffff" after 47.823911955977984us,
    X"ffffffff" after 47.92396198099049us,
    X"ffffffff" after 48.024012006003us,
    X"ffffffff" after 48.124062031015505us,
    X"ffffffff" after 48.22411205602801us,
    X"ffffffff" after 48.32416208104052us,
    X"ffffffff" after 48.42421210605303us,
    X"ffffffff" after 48.52426213106553us,
    X"ffffffff" after 48.624312156078034us,
    X"ffffffff" after 48.72436218109054us,
    X"ffffffff" after 48.82441220610305us,
    X"ffffffff" after 48.924462231115555us,
    X"ffffffff" after 49.02451225612806us,
    X"ffffffff" after 49.12456228114057us,
    X"ffffffff" after 49.22461230615308us,
    X"ffffffff" after 49.32466233116558us,
    X"ffffffff" after 49.424712356178084us,
    X"ffffffff" after 49.52476238119059us,
    X"ffffffff" after 49.6248124062031us,
    X"ffffffff" after 49.724862431215605us,
    X"ffffffff" after 49.82491245622811us,
    X"ffffffff" after 49.92496248124062us,
    X"ffffffff" after 50.02501250625313us,
    X"ffffffff" after 50.12506253126563us,
    X"ffffffff" after 50.225112556278134us,
    X"ffffffff" after 50.32516258129064us,
    X"ffffffff" after 50.42521260630315us,
    X"ffffffff" after 50.525262631315655us,
    X"ffffffff" after 50.62531265632816us,
    X"ffffffff" after 50.72536268134067us,
    X"ffffffff" after 50.82541270635318us,
    X"ffffffff" after 50.92546273136568us,
    X"ffffffff" after 51.025512756378184us,
    X"ffffffff" after 51.12556278139069us,
    X"ffffffff" after 51.2256128064032us,
    X"ffffffff" after 51.325662831415706us,
    X"ffffffff" after 51.42571285642821us,
    X"ffffffff" after 51.52576288144072us,
    X"ffffffff" after 51.62581290645322us,
    X"ffffffff" after 51.72586293146573us,
    X"ffffffff" after 51.825912956478234us,
    X"ffffffff" after 51.92596298149074us,
    X"ffffffff" after 52.02601300650325us,
    X"ffffffff" after 52.126063031515756us,
    X"ffffffff" after 52.22611305652826us,
    X"ffffffff" after 52.32616308154077us,
    X"ffffffff" after 52.42621310655327us,
    X"ffffffff" after 52.52626313156578us,
    X"ffffffff" after 52.626313156578284us,
    X"ffffffff" after 52.72636318159079us,
    X"ffffffff" after 52.8264132066033us,
    X"ffffffff" after 52.926463231615806us,
    X"ffffffff" after 53.02651325662831us,
    X"ffffffff" after 53.12656328164082us,
    X"ffffffff" after 53.22661330665332us,
    X"ffffffff" after 53.32666333166583us,
    X"ffffffff" after 53.426713356678334us,
    X"ffffffff" after 53.52676338169084us,
    X"ffffffff" after 53.62681340670335us,
    X"ffffffff" after 53.726863431715856us,
    X"ffffffff" after 53.82691345672836us,
    X"ffffffff" after 53.92696348174087us,
    X"ffffffff" after 54.02701350675337us,
    X"ffffffff" after 54.12706353176588us,
    X"ffffffff" after 54.227113556778384us,
    X"ffffffff" after 54.32716358179089us,
    X"ffffffff" after 54.4272136068034us,
    X"ffffffff" after 54.527263631815906us,
    X"ffffffff" after 54.62731365682841us,
    X"ffffffff" after 54.72736368184092us,
    X"ffffffff" after 54.82741370685342us,
    X"ffffffff" after 54.92746373186593us,
    X"ffffffff" after 55.027513756878434us,
    X"ffffffff" after 55.12756378189094us,
    X"ffffffff" after 55.22761380690345us,
    X"ffffffff" after 55.327663831915956us,
    X"ffffffff" after 55.42771385692846us,
    X"ffffffff" after 55.52776388194097us,
    X"ffffffff" after 55.62781390695347us,
    X"ffffffff" after 55.72786393196598us,
    X"ffffffff" after 55.827913956978485us,
    X"ffffffff" after 55.92796398199099us,
    X"ffffffff" after 56.0280140070035us,
    X"ffffffff" after 56.128064032016006us,
    X"ffffffff" after 56.22811405702851us,
    X"ffffffff" after 56.32816408204102us,
    X"ffffffff" after 56.42821410705352us,
    X"ffffffff" after 56.52826413206603us,
    X"ffffffff" after 56.628314157078535us,
    X"ffffffff" after 56.72836418209104us,
    X"ffffffff" after 56.82841420710355us,
    X"ffffffff" after 56.928464232116056us,
    X"ffffffff" after 57.02851425712856us,
    X"ffffffff" after 57.12856428214107us,
    X"ffffffff" after 57.22861430715357us,
    X"ffffffff" after 57.32866433216608us,
    X"ffffffff" after 57.428714357178585us,
    X"ffffffff" after 57.52876438219109us,
    X"ffffffff" after 57.6288144072036us,
    X"ffffffff" after 57.728864432216106us,
    X"ffffffff" after 57.82891445722861us,
    X"ffffffff" after 57.92896448224111us,
    X"ffffffff" after 58.02901450725362us,
    X"ffffffff" after 58.12906453226613us,
    X"ffffffff" after 58.229114557278635us,
    X"ffffffff" after 58.32916458229114us,
    X"ffffffff" after 58.42921460730365us,
    X"ffffffff" after 58.529264632316156us,
    X"ffffffff" after 58.62931465732866us,
    X"ffffffff" after 58.72936468234116us,
    X"ffffffff" after 58.82941470735367us,
    X"ffffffff" after 58.92946473236618us,
    X"ffffffff" after 59.029514757378685us,
    X"ffffffff" after 59.12956478239119us,
    X"ffffffff" after 59.2296148074037us,
    X"ffffffff" after 59.329664832416206us,
    X"ffffffff" after 59.42971485742871us,
    X"ffffffff" after 59.529764882441214us,
    X"ffffffff" after 59.62981490745372us,
    X"ffffffff" after 59.72986493246623us,
    X"ffffffff" after 59.829914957478735us,
    X"ffffffff" after 59.92996498249124us,
    X"ffffffff" after 60.03001500750375us,
    X"ffffffff" after 60.13006503251626us,
    X"ffffffff" after 60.230115057528764us,
    X"ffffffff" after 60.330165082541264us,
    X"ffffffff" after 60.43021510755377us,
    X"ffffffff" after 60.53026513256628us,
    X"ffffffff" after 60.630315157578785us,
    X"ffffffff" after 60.73036518259129us,
    X"ffffffff" after 60.8304152076038us,
    X"ffffffff" after 60.93046523261631us,
    X"ffffffff" after 61.030515257628814us,
    X"ffffffff" after 61.130565282641314us,
    X"ffffffff" after 61.23061530765382us,
    X"ffffffff" after 61.33066533266633us,
    X"ffffffff" after 61.430715357678835us,
    X"ffffffff" after 61.53076538269134us,
    X"ffffffff" after 61.63081540770385us,
    X"ffffffff" after 61.73086543271636us,
    X"ffffffff" after 61.830915457728864us,
    X"ffffffff" after 61.930965482741364us,
    X"ffffffff" after 62.03101550775387us,
    X"ffffffff" after 62.13106553276638us,
    X"ffffffff" after 62.231115557778885us,
    X"ffffffff" after 62.33116558279139us,
    X"ffffffff" after 62.4312156078039us,
    X"ffffffff" after 62.53126563281641us,
    X"ffffffff" after 62.631315657828914us,
    X"ffffffff" after 62.731365682841414us,
    X"ffffffff" after 62.83141570785392us,
    X"ffffffff" after 62.93146573286643us,
    X"ffffffff" after 63.031515757878935us,
    X"ffffffff" after 63.13156578289144us,
    X"ffffffff" after 63.23161580790395us,
    X"ffffffff" after 63.33166583291646us,
    X"ffffffff" after 63.431715857928964us,
    X"ffffffff" after 63.531765882941464us,
    X"ffffffff" after 63.63181590795397us,
    X"ffffffff" after 63.73186593296648us,
    X"ffffffff" after 63.831915957978985us,
    X"ffffffff" after 63.93196598299149us,
    X"ffffffff" after 64.03201600800399us,
    X"ffffffff" after 64.1320660330165us,
    X"ffffffff" after 64.232116058029us,
    X"ffffffff" after 64.33216608304151us,
    X"ffffffff" after 64.43221610805402us,
    X"ffffffff" after 64.53226613306653us,
    X"ffffffff" after 64.63231615807904us,
    X"ffffffff" after 64.73236618309154us,
    X"ffffffff" after 64.83241620810405us,
    X"ffffffff" after 64.93246623311656us,
    X"ffffffff" after 65.03251625812906us,
    X"ffffffff" after 65.13256628314157us,
    X"ffffffff" after 65.23261630815408us,
    X"ffffffff" after 65.33266633316659us,
    X"ffffffff" after 65.43271635817908us,
    X"ffffffff" after 65.53276638319159us,
    X"ffffffff" after 65.63281640820409us,
    X"ffffffff" after 65.7328664332166us,
    X"ffffffff" after 65.8329164582291us,
    X"ffffffff" after 65.93296648324161us,
    X"ffffffff" after 66.03301650825412us,
    X"ffffffff" after 66.13306653326663us,
    X"ffffffff" after 66.23311655827914us,
    X"ffffffff" after 66.33316658329164us,
    X"ffffffff" after 66.43321660830415us,
    X"ffffffff" after 66.53326663331666us,
    X"ffffffff" after 66.63331665832916us,
    X"ffffffff" after 66.73336668334167us,
    X"ffffffff" after 66.83341670835418us,
    X"ffffffff" after 66.93346673336669us,
    X"ffffffff" after 67.03351675837918us,
    X"ffffffff" after 67.13356678339169us,
    X"ffffffff" after 67.2336168084042us,
    X"ffffffff" after 67.3336668334167us,
    X"ffffffff" after 67.43371685842921us,
    X"ffffffff" after 67.53376688344171us,
    X"ffffffff" after 67.63381690845422us,
    X"ffffffff" after 67.73386693346673us,
    X"ffffffff" after 67.83391695847924us,
    X"ffffffff" after 67.93396698349174us,
    X"ffffffff" after 68.03401700850425us,
    X"ffffffff" after 68.13406703351676us,
    X"ffffffff" after 68.23411705852926us,
    X"ffffffff" after 68.33416708354177us,
    X"ffffffff" after 68.43421710855428us,
    X"ffffffff" after 68.53426713356679us,
    X"ffffffff" after 68.63431715857928us,
    X"ffffffff" after 68.73436718359179us,
    X"ffffffff" after 68.8344172086043us,
    X"ffffffff" after 68.9344672336168us,
    X"ffffffff" after 69.03451725862931us,
    X"ffffffff" after 69.13456728364181us,
    X"ffffffff" after 69.23461730865432us,
    X"ffffffff" after 69.33466733366683us,
    X"ffffffff" after 69.43471735867934us,
    X"ffffffff" after 69.53476738369184us,
    X"ffffffff" after 69.63481740870435us,
    X"ffffffff" after 69.73486743371686us,
    X"ffffffff" after 69.83491745872936us,
    X"ffffffff" after 69.93496748374187us,
    X"ffffffff" after 70.03501750875438us,
    X"ffffffff" after 70.13506753376689us,
    X"ffffffff" after 70.23511755877938us,
    X"ffffffff" after 70.33516758379189us,
    X"ffffffff" after 70.4352176088044us,
    X"ffffffff" after 70.5352676338169us,
    X"ffffffff" after 70.63531765882941us,
    X"ffffffff" after 70.73536768384191us,
    X"ffffffff" after 70.83541770885442us,
    X"ffffffff" after 70.93546773386693us,
    X"ffffffff" after 71.03551775887944us,
    X"ffffffff" after 71.13556778389194us,
    X"ffffffff" after 71.23561780890445us,
    X"ffffffff" after 71.33566783391696us,
    X"ffffffff" after 71.43571785892946us,
    X"ffffffff" after 71.53576788394197us,
    X"ffffffff" after 71.63581790895448us,
    X"ffffffff" after 71.73586793396697us,
    X"ffffffff" after 71.83591795897948us,
    X"ffffffff" after 71.93596798399199us,
    X"ffffffff" after 72.0360180090045us,
    X"ffffffff" after 72.136068034017us,
    X"ffffffff" after 72.23611805902951us,
    X"ffffffff" after 72.33616808404201us,
    X"ffffffff" after 72.43621810905452us,
    X"ffffffff" after 72.53626813406703us,
    X"ffffffff" after 72.63631815907954us,
    X"ffffffff" after 72.73636818409204us,
    X"ffffffff" after 72.83641820910455us,
    X"ffffffff" after 72.93646823411706us,
    X"ffffffff" after 73.03651825912956us,
    X"ffffffff" after 73.13656828414207us,
    X"ffffffff" after 73.23661830915458us,
    X"ffffffff" after 73.33666833416707us,
    X"ffffffff" after 73.43671835917958us,
    X"ffffffff" after 73.53676838419209us,
    X"ffffffff" after 73.6368184092046us,
    X"ffffffff" after 73.7368684342171us,
    X"ffffffff" after 73.83691845922961us,
    X"ffffffff" after 73.93696848424212us,
    X"ffffffff" after 74.03701850925462us,
    X"ffffffff" after 74.13706853426713us,
    X"ffffffff" after 74.23711855927964us,
    X"ffffffff" after 74.33716858429214us,
    X"ffffffff" after 74.43721860930465us,
    X"ffffffff" after 74.53726863431716us,
    X"ffffffff" after 74.63731865932967us,
    X"ffffffff" after 74.73736868434217us,
    X"ffffffff" after 74.83741870935468us,
    X"ffffffff" after 74.93746873436717us,
    X"ffffffff" after 75.03751875937968us,
    X"ffffffff" after 75.13756878439219us,
    X"ffffffff" after 75.2376188094047us,
    X"ffffffff" after 75.3376688344172us,
    X"ffffffff" after 75.43771885942971us,
    X"ffffffff" after 75.53776888444222us,
    X"ffffffff" after 75.63781890945472us,
    X"ffffffff" after 75.73786893446723us,
    X"ffffffff" after 75.83791895947974us,
    X"ffffffff" after 75.93796898449224us,
    X"ffffffff" after 76.03801900950475us,
    X"ffffffff" after 76.13806903451726us,
    X"ffffffff" after 76.23811905952977us,
    X"ffffffff" after 76.33816908454227us,
    X"ffffffff" after 76.43821910955478us,
    X"ffffffff" after 76.53826913456727us,
    X"ffffffff" after 76.63831915957978us,
    X"ffffffff" after 76.73836918459229us,
    X"ffffffff" after 76.8384192096048us,
    X"ffffffff" after 76.9384692346173us,
    X"ffffffff" after 77.03851925962981us,
    X"ffffffff" after 77.13856928464232us,
    X"ffffffff" after 77.23861930965482us,
    X"ffffffff" after 77.33866933466733us,
    X"ffffffff" after 77.43871935967984us,
    X"ffffffff" after 77.53876938469234us,
    X"ffffffff" after 77.63881940970485us,
    X"ffffffff" after 77.73886943471736us,
    X"ffffffff" after 77.83891945972987us,
    X"ffffffff" after 77.93896948474237us,
    X"ffffffff" after 78.03901950975487us,
    X"ffffffff" after 78.13906953476737us,
    X"ffffffff" after 78.23911955977988us,
    X"ffffffff" after 78.33916958479239us,
    X"ffffffff" after 78.4392196098049us,
    X"ffffffff" after 78.5392696348174us,
    X"ffffffff" after 78.63931965982991us,
    X"ffffffff" after 78.73936968484242us,
    X"ffffffff" after 78.83941970985492us,
    X"ffffffff" after 78.93946973486743us,
    X"ffffffff" after 79.03951975987994us,
    X"ffffffff" after 79.13956978489244us,
    X"ffffffff" after 79.23961980990495us,
    X"ffffffff" after 79.33966983491746us,
    X"ffffffff" after 79.43971985992997us,
    X"ffffffff" after 79.53976988494247us,
    X"ffffffff" after 79.63981990995497us,
    X"ffffffff" after 79.73986993496747us,
    X"ffffffff" after 79.83991995997998us,
    X"ffffffff" after 79.93996998499249us,
    X"ffffffff" after 80.040020010005us,
    X"ffffffff" after 80.1400700350175us,
    X"ffffffff" after 80.24012006003001us,
    X"ffffffff" after 80.34017008504252us,
    X"ffffffff" after 80.44022011005502us,
    X"ffffffff" after 80.54027013506753us,
    X"ffffffff" after 80.64032016008004us,
    X"ffffffff" after 80.74037018509254us,
    X"ffffffff" after 80.84042021010505us,
    X"ffffffff" after 80.94047023511756us,
    X"ffffffff" after 81.04052026013007us,
    X"ffffffff" after 81.14057028514257us,
    X"ffffffff" after 81.24062031015507us,
    X"ffffffff" after 81.34067033516757us,
    X"ffffffff" after 81.44072036018008us,
    X"ffffffff" after 81.54077038519259us,
    X"ffffffff" after 81.6408204102051us,
    X"ffffffff" after 81.7408704352176us,
    X"ffffffff" after 81.84092046023011us,
    X"ffffffff" after 81.94097048524262us,
    X"ffffffff" after 82.04102051025512us,
    X"ffffffff" after 82.14107053526763us,
    X"ffffffff" after 82.24112056028014us,
    X"ffffffff" after 82.34117058529264us,
    X"ffffffff" after 82.44122061030515us,
    X"ffffffff" after 82.54127063531766us,
    X"ffffffff" after 82.64132066033017us,
    X"ffffffff" after 82.74137068534267us,
    X"ffffffff" after 82.84142071035517us,
    X"ffffffff" after 82.94147073536767us,
    X"ffffffff" after 83.04152076038018us,
    X"ffffffff" after 83.14157078539269us,
    X"ffffffff" after 83.2416208104052us,
    X"ffffffff" after 83.3416708354177us,
    X"ffffffff" after 83.44172086043021us,
    X"ffffffff" after 83.54177088544272us,
    X"ffffffff" after 83.64182091045522us,
    X"ffffffff" after 83.74187093546773us,
    X"ffffffff" after 83.84192096048024us,
    X"ffffffff" after 83.94197098549274us,
    X"ffffffff" after 84.04202101050525us,
    X"ffffffff" after 84.14207103551776us,
    X"ffffffff" after 84.24212106053027us,
    X"ffffffff" after 84.34217108554276us,
    X"ffffffff" after 84.44222111055527us,
    X"ffffffff" after 84.54227113556777us,
    X"ffffffff" after 84.64232116058028us,
    X"ffffffff" after 84.74237118559279us,
    X"ffffffff" after 84.8424212106053us,
    X"ffffffff" after 84.9424712356178us,
    X"ffffffff" after 85.04252126063031us,
    X"ffffffff" after 85.14257128564282us,
    X"ffffffff" after 85.24262131065532us,
    X"ffffffff" after 85.34267133566783us,
    X"ffffffff" after 85.44272136068034us,
    X"ffffffff" after 85.54277138569284us,
    X"ffffffff" after 85.64282141070535us,
    X"ffffffff" after 85.74287143571786us,
    X"ffffffff" after 85.84292146073037us,
    X"ffffffff" after 85.94297148574286us,
    X"ffffffff" after 86.04302151075537us,
    X"ffffffff" after 86.14307153576787us,
    X"ffffffff" after 86.24312156078038us,
    X"ffffffff" after 86.34317158579289us,
    X"ffffffff" after 86.4432216108054us,
    X"ffffffff" after 86.5432716358179us,
    X"ffffffff" after 86.64332166083041us,
    X"ffffffff" after 86.74337168584292us,
    X"ffffffff" after 86.84342171085542us,
    X"ffffffff" after 86.94347173586793us,
    X"ffffffff" after 87.04352176088044us,
    X"ffffffff" after 87.14357178589295us,
    X"ffffffff" after 87.24362181090545us,
    X"ffffffff" after 87.34367183591796us,
    X"ffffffff" after 87.44372186093047us,
    X"ffffffff" after 87.54377188594296us,
    X"ffffffff" after 87.64382191095547us,
    X"ffffffff" after 87.74387193596797us,
    X"ffffffff" after 87.84392196098048us,
    X"ffffffff" after 87.94397198599299us,
    X"ffffffff" after 88.0440220110055us,
    X"ffffffff" after 88.144072036018us,
    X"ffffffff" after 88.24412206103051us,
    X"ffffffff" after 88.34417208604302us,
    X"ffffffff" after 88.44422211105552us,
    X"ffffffff" after 88.54427213606803us,
    X"ffffffff" after 88.64432216108054us,
    X"ffffffff" after 88.74437218609305us,
    X"ffffffff" after 88.84442221110555us,
    X"ffffffff" after 88.94447223611806us,
    X"ffffffff" after 89.04452226113057us,
    X"ffffffff" after 89.14457228614306us,
    X"ffffffff" after 89.24462231115557us,
    X"ffffffff" after 89.34467233616807us,
    X"ffffffff" after 89.44472236118058us,
    X"ffffffff" after 89.54477238619309us,
    X"ffffffff" after 89.6448224112056us,
    X"ffffffff" after 89.7448724362181us,
    X"ffffffff" after 89.84492246123061us,
    X"ffffffff" after 89.94497248624312us,
    X"ffffffff" after 90.04502251125562us,
    X"ffffffff" after 90.14507253626813us,
    X"ffffffff" after 90.24512256128064us,
    X"ffffffff" after 90.34517258629315us,
    X"ffffffff" after 90.44522261130565us,
    X"ffffffff" after 90.54527263631816us,
    X"ffffffff" after 90.64532266133065us,
    X"ffffffff" after 90.74537268634316us,
    X"ffffffff" after 90.84542271135567us,
    X"ffffffff" after 90.94547273636817us,
    X"ffffffff" after 91.04552276138068us,
    X"ffffffff" after 91.14557278639319us,
    X"ffffffff" after 91.2456228114057us,
    X"ffffffff" after 91.3456728364182us,
    X"ffffffff" after 91.44572286143071us,
    X"ffffffff" after 91.54577288644322us,
    X"ffffffff" after 91.64582291145572us,
    X"ffffffff" after 91.74587293646823us,
    X"ffffffff" after 91.84592296148074us,
    X"ffffffff" after 91.94597298649325us,
    X"ffffffff" after 92.04602301150575us,
    X"ffffffff" after 92.14607303651826us,
    X"ffffffff" after 92.24612306153075us,
    X"ffffffff" after 92.34617308654326us,
    X"ffffffff" after 92.44622311155577us,
    X"ffffffff" after 92.54627313656827us,
    X"ffffffff" after 92.64632316158078us,
    X"ffffffff" after 92.74637318659329us,
    X"ffffffff" after 92.8464232116058us,
    X"ffffffff" after 92.9464732366183us,
    X"ffffffff" after 93.04652326163081us,
    X"ffffffff" after 93.14657328664332us,
    X"ffffffff" after 93.24662331165582us,
    X"ffffffff" after 93.34667333666833us,
    X"ffffffff" after 93.44672336168084us,
    X"ffffffff" after 93.54677338669335us,
    X"ffffffff" after 93.64682341170585us,
    X"ffffffff" after 93.74687343671836us,
    X"ffffffff" after 93.84692346173085us,
    X"ffffffff" after 93.94697348674336us,
    X"ffffffff" after 94.04702351175587us,
    X"ffffffff" after 94.14707353676837us,
    X"ffffffff" after 94.24712356178088us,
    X"ffffffff" after 94.34717358679339us,
    X"ffffffff" after 94.4472236118059us,
    X"ffffffff" after 94.5472736368184us,
    X"ffffffff" after 94.64732366183091us,
    X"ffffffff" after 94.74737368684342us,
    X"ffffffff" after 94.84742371185592us,
    X"ffffffff" after 94.94747373686843us,
    X"ffffffff" after 95.04752376188094us,
    X"ffffffff" after 95.14757378689345us,
    X"ffffffff" after 95.24762381190595us,
    X"ffffffff" after 95.34767383691846us,
    X"ffffffff" after 95.44772386193095us,
    X"ffffffff" after 95.54777388694346us,
    X"ffffffff" after 95.64782391195597us,
    X"ffffffff" after 95.74787393696847us,
    X"ffffffff" after 95.84792396198098us,
    X"ffffffff" after 95.94797398699349us,
    X"ffffffff" after 96.048024012006us,
    X"ffffffff" after 96.1480740370185us,
    X"ffffffff" after 96.24812406203101us,
    X"ffffffff" after 96.34817408704352us,
    X"ffffffff" after 96.44822411205602us,
    X"ffffffff" after 96.54827413706853us,
    X"ffffffff" after 96.64832416208104us,
    X"ffffffff" after 96.74837418709355us,
    X"ffffffff" after 96.84842421210605us,
    X"ffffffff" after 96.94847423711855us,
    X"ffffffff" after 97.04852426213105us,
    X"ffffffff" after 97.14857428714356us,
    X"ffffffff" after 97.24862431215607us,
    X"ffffffff" after 97.34867433716857us,
    X"ffffffff" after 97.44872436218108us,
    X"ffffffff" after 97.54877438719359us,
    X"ffffffff" after 97.6488244122061us,
    X"ffffffff" after 97.7488744372186us,
    X"ffffffff" after 97.84892446223111us,
    X"ffffffff" after 97.94897448724362us,
    X"ffffffff" after 98.04902451225612us,
    X"ffffffff" after 98.14907453726863us,
    X"ffffffff" after 98.24912456228114us,
    X"ffffffff" after 98.34917458729365us,
    X"ffffffff" after 98.44922461230615us,
    X"ffffffff" after 98.54927463731865us,
    X"ffffffff" after 98.64932466233115us,
    X"ffffffff" after 98.74937468734366us,
    X"ffffffff" after 98.84942471235617us,
    X"ffffffff" after 98.94947473736867us,
    X"ffffffff" after 99.04952476238118us,
    X"ffffffff" after 99.14957478739369us,
    X"ffffffff" after 99.2496248124062us,
    X"ffffffff" after 99.3496748374187us,
    X"ffffffff" after 99.44972486243121us,
    X"ffffffff" after 99.54977488744372us,
    X"ffffffff" after 99.64982491245622us,
    X"ffffffff" after 99.74987493746873us,
    X"ffffffff" after 99.84992496248124us,
    X"ffffffff" after 99.94997498749375us,
    X"7f800000" after 100.05002501250625us,
    X"7f800000" after 100.15007503751875us,
    X"7f800000" after 100.25012506253125us,
    X"7f800000" after 100.35017508754376us,
    X"7f800000" after 100.45022511255627us,
    X"7f800000" after 100.55027513756878us,
    X"7f800000" after 100.65032516258128us,
    X"7f800000" after 100.75037518759379us,
    X"7f800000" after 100.8504252126063us,
    X"7f800000" after 100.9504752376188us,
    X"7f800000" after 101.05052526263131us,
    X"7f800000" after 101.15057528764382us,
    X"7f800000" after 101.25062531265633us,
    X"7f800000" after 101.35067533766883us,
    X"7f800000" after 101.45072536268134us,
    X"7f800000" after 101.55077538769385us,
    X"7f800000" after 101.65082541270635us,
    X"7f800000" after 101.75087543771885us,
    X"7f800000" after 101.85092546273135us,
    X"7f800000" after 101.95097548774386us,
    X"7f800000" after 102.05102551275637us,
    X"7f800000" after 102.15107553776888us,
    X"7f800000" after 102.25112556278138us,
    X"7f800000" after 102.35117558779389us,
    X"7f800000" after 102.4512256128064us,
    X"7f800000" after 102.5512756378189us,
    X"7f800000" after 102.65132566283141us,
    X"7f800000" after 102.75137568784392us,
    X"7f800000" after 102.85142571285643us,
    X"7f800000" after 102.95147573786893us,
    X"7f800000" after 103.05152576288144us,
    X"7f800000" after 103.15157578789395us,
    X"7f800000" after 103.25162581290644us,
    X"7f800000" after 103.35167583791895us,
    X"7f800000" after 103.45172586293145us,
    X"7f800000" after 103.55177588794396us,
    X"7f800000" after 103.65182591295647us,
    X"7f800000" after 103.75187593796898us,
    X"7f800000" after 103.85192596298148us,
    X"7f800000" after 103.95197598799399us,
    X"7f800000" after 104.0520260130065us,
    X"7f800000" after 104.152076038019us,
    X"7f800000" after 104.25212606303151us,
    X"7f800000" after 104.35217608804402us,
    X"7f800000" after 104.45222611305653us,
    X"7f800000" after 104.55227613806903us,
    X"7f800000" after 104.65232616308154us,
    X"7f800000" after 104.75237618809405us,
    X"7f800000" after 104.85242621310654us,
    X"7f800000" after 104.95247623811905us,
    X"7f800000" after 105.05252626313155us,
    X"7f800000" after 105.15257628814406us,
    X"7f800000" after 105.25262631315657us,
    X"7f800000" after 105.35267633816908us,
    X"7f800000" after 105.45272636318158us,
    X"7f800000" after 105.55277638819409us,
    X"7f800000" after 105.6528264132066us,
    X"7f800000" after 105.7528764382191us,
    X"7f800000" after 105.85292646323161us,
    X"7f800000" after 105.95297648824412us,
    X"7f800000" after 106.05302651325663us,
    X"7f800000" after 106.15307653826913us,
    X"7f800000" after 106.25312656328164us,
    X"7f800000" after 106.35317658829415us,
    X"7f800000" after 106.45322661330664us,
    X"7f800000" after 106.55327663831915us,
    X"7f800000" after 106.65332666333165us,
    X"7f800000" after 106.75337668834416us,
    X"7f800000" after 106.85342671335667us,
    X"7f800000" after 106.95347673836918us,
    X"7f800000" after 107.05352676338168us,
    X"7f800000" after 107.15357678839419us,
    X"7f800000" after 107.2536268134067us,
    X"7f800000" after 107.3536768384192us,
    X"7f800000" after 107.45372686343171us,
    X"7f800000" after 107.55377688844422us,
    X"7f800000" after 107.65382691345673us,
    X"7f800000" after 107.75387693846923us,
    X"7f800000" after 107.85392696348174us,
    X"7f800000" after 107.95397698849425us,
    X"7f800000" after 108.05402701350674us,
    X"7f800000" after 108.15407703851925us,
    X"7f800000" after 108.25412706353175us,
    X"7f800000" after 108.35417708854426us,
    X"7f800000" after 108.45422711355677us,
    X"7f800000" after 108.55427713856928us,
    X"7f800000" after 108.65432716358178us,
    X"7f800000" after 108.75437718859429us,
    X"7f800000" after 108.8544272136068us,
    X"7f800000" after 108.9544772386193us,
    X"7f800000" after 109.05452726363181us,
    X"7f800000" after 109.15457728864432us,
    X"7f800000" after 109.25462731365683us,
    X"7f800000" after 109.35467733866933us,
    X"7f800000" after 109.45472736368184us,
    X"7f800000" after 109.55477738869433us,
    X"7f800000" after 109.65482741370684us,
    X"7f800000" after 109.75487743871935us,
    X"7f800000" after 109.85492746373185us,
    X"7f800000" after 109.95497748874436us,
    X"ffffffff" after 110.05502751375687us,
    X"ffffffff" after 110.15507753876938us,
    X"ffffffff" after 110.25512756378188us,
    X"ffffffff" after 110.35517758879439us,
    X"ffffffff" after 110.4552276138069us,
    X"ffffffff" after 110.5552776388194us,
    X"ffffffff" after 110.65532766383191us,
    X"ffffffff" after 110.75537768884442us,
    X"ffffffff" after 110.85542771385693us,
    X"ffffffff" after 110.95547773886943us,
    X"ffffffff" after 111.05552776388194us,
    X"ffffffff" after 111.15557778889443us,
    X"ffffffff" after 111.25562781390694us,
    X"ffffffff" after 111.35567783891945us,
    X"ffffffff" after 111.45572786393195us,
    X"ffffffff" after 111.55577788894446us,
    X"ffffffff" after 111.65582791395697us,
    X"ffffffff" after 111.75587793896948us,
    X"ffffffff" after 111.85592796398198us,
    X"ffffffff" after 111.95597798899449us,
    X"ffffffff" after 112.056028014007us,
    X"ffffffff" after 112.1560780390195us,
    X"ffffffff" after 112.25612806403201us,
    X"ffffffff" after 112.35617808904452us,
    X"ffffffff" after 112.45622811405703us,
    X"ffffffff" after 112.55627813906953us,
    X"ffffffff" after 112.65632816408204us,
    X"ffffffff" after 112.75637818909453us,
    X"ffffffff" after 112.85642821410704us,
    X"ffffffff" after 112.95647823911955us,
    X"ffffffff" after 113.05652826413206us,
    X"ffffffff" after 113.15657828914456us,
    X"ffffffff" after 113.25662831415707us,
    X"ffffffff" after 113.35667833916958us,
    X"ffffffff" after 113.45672836418208us,
    X"ffffffff" after 113.55677838919459us,
    X"ffffffff" after 113.6568284142071us,
    X"ffffffff" after 113.7568784392196us,
    X"ffffffff" after 113.85692846423211us,
    X"ffffffff" after 113.95697848924462us,
    X"ffffffff" after 114.05702851425713us,
    X"ffffffff" after 114.15707853926963us,
    X"ffffffff" after 114.25712856428214us,
    X"ffffffff" after 114.35717858929463us,
    X"ffffffff" after 114.45722861430714us,
    X"ffffffff" after 114.55727863931965us,
    X"ffffffff" after 114.65732866433216us,
    X"ffffffff" after 114.75737868934466us,
    X"ffffffff" after 114.85742871435717us,
    X"ffffffff" after 114.95747873936968us,
    X"ffffffff" after 115.05752876438218us,
    X"ffffffff" after 115.15757878939469us,
    X"ffffffff" after 115.2576288144072us,
    X"ffffffff" after 115.3576788394197us,
    X"ffffffff" after 115.45772886443221us,
    X"ffffffff" after 115.55777888944472us,
    X"ffffffff" after 115.65782891445723us,
    X"ffffffff" after 115.75787893946973us,
    X"ffffffff" after 115.85792896448223us,
    X"ffffffff" after 115.95797898949473us,
    X"ffffffff" after 116.05802901450724us,
    X"ffffffff" after 116.15807903951975us,
    X"ffffffff" after 116.25812906453226us,
    X"ffffffff" after 116.35817908954476us,
    X"ffffffff" after 116.45822911455727us,
    X"ffffffff" after 116.55827913956978us,
    X"ffffffff" after 116.65832916458228us,
    X"ffffffff" after 116.75837918959479us,
    X"ffffffff" after 116.8584292146073us,
    X"ffffffff" after 116.9584792396198us,
    X"ffffffff" after 117.05852926463231us,
    X"ffffffff" after 117.15857928964482us,
    X"ffffffff" after 117.25862931465733us,
    X"ffffffff" after 117.35867933966983us,
    X"ffffffff" after 117.45872936468233us,
    X"ffffffff" after 117.55877938969483us,
    X"ffffffff" after 117.65882941470734us,
    X"ffffffff" after 117.75887943971985us,
    X"ffffffff" after 117.85892946473236us,
    X"ffffffff" after 117.95897948974486us,
    X"ffffffff" after 118.05902951475737us,
    X"ffffffff" after 118.15907953976988us,
    X"ffffffff" after 118.25912956478238us,
    X"ffffffff" after 118.35917958979489us,
    X"ffffffff" after 118.4592296148074us,
    X"ffffffff" after 118.5592796398199us,
    X"ffffffff" after 118.65932966483241us,
    X"ffffffff" after 118.75937968984492us,
    X"ffffffff" after 118.85942971485743us,
    X"ffffffff" after 118.95947973986993us,
    X"ffffffff" after 119.05952976488243us,
    X"ffffffff" after 119.15957978989493us,
    X"ffffffff" after 119.25962981490744us,
    X"ffffffff" after 119.35967983991995us,
    X"ffffffff" after 119.45972986493246us,
    X"ffffffff" after 119.55977988994496us,
    X"ffffffff" after 119.65982991495747us,
    X"ffffffff" after 119.75987993996998us,
    X"ffffffff" after 119.85992996498248us,
    X"ffffffff" after 119.95997998999499us,
    X"ffffffff" after 120.0600300150075us,
    X"ffffffff" after 120.16008004002us,
    X"ffffffff" after 120.26013006503251us,
    X"ffffffff" after 120.36018009004502us,
    X"ffffffff" after 120.46023011505753us,
    X"ffffffff" after 120.56028014007003us,
    X"ffffffff" after 120.66033016508253us,
    X"ffffffff" after 120.76038019009503us,
    X"ffffffff" after 120.86043021510754us,
    X"ffffffff" after 120.96048024012005us,
    X"ffffffff" after 121.06053026513256us,
    X"ffffffff" after 121.16058029014506us,
    X"ffffffff" after 121.26063031515757us,
    X"ffffffff" after 121.36068034017008us,
    X"ffffffff" after 121.46073036518258us,
    X"ffffffff" after 121.56078039019509us,
    X"ffffffff" after 121.6608304152076us,
    X"ffffffff" after 121.7608804402201us,
    X"ffffffff" after 121.86093046523261us,
    X"ffffffff" after 121.96098049024512us,
    X"ffffffff" after 122.06103051525763us,
    X"ffffffff" after 122.16108054027012us,
    X"ffffffff" after 122.26113056528263us,
    X"ffffffff" after 122.36118059029513us,
    X"ffffffff" after 122.46123061530764us,
    X"ffffffff" after 122.56128064032015us,
    X"ffffffff" after 122.66133066533266us,
    X"ffffffff" after 122.76138069034516us,
    X"ffffffff" after 122.86143071535767us,
    X"ffffffff" after 122.96148074037018us,
    X"ffffffff" after 123.06153076538268us,
    X"ffffffff" after 123.16158079039519us,
    X"ffffffff" after 123.2616308154077us,
    X"ffffffff" after 123.3616808404202us,
    X"ffffffff" after 123.46173086543271us,
    X"ffffffff" after 123.56178089044522us,
    X"ffffffff" after 123.66183091545773us,
    X"ffffffff" after 123.76188094047022us,
    X"ffffffff" after 123.86193096548273us,
    X"ffffffff" after 123.96198099049523us,
    X"ffffffff" after 124.06203101550774us,
    X"ffffffff" after 124.16208104052025us,
    X"ffffffff" after 124.26213106553276us,
    X"ffffffff" after 124.36218109054526us,
    X"ffffffff" after 124.46223111555777us,
    X"ffffffff" after 124.56228114057028us,
    X"ffffffff" after 124.66233116558278us,
    X"ffffffff" after 124.76238119059529us,
    X"ffffffff" after 124.8624312156078us,
    X"ffffffff" after 124.9624812406203us,
    X"26400000" after 125.06253126563281us,
    X"26400000" after 125.16258129064532us,
    X"26400000" after 125.26263131565783us,
    X"26400000" after 125.36268134067032us,
    X"26400000" after 125.46273136568283us,
    X"26400000" after 125.56278139069533us,
    X"26400000" after 125.66283141570784us,
    X"26400000" after 125.76288144072035us,
    X"26400000" after 125.86293146573286us,
    X"26400000" after 125.96298149074536us,
    X"26400000" after 126.06303151575787us,
    X"26400000" after 126.16308154077038us,
    X"26400000" after 126.26313156578288us,
    X"26400000" after 126.36318159079539us,
    X"26400000" after 126.4632316158079us,
    X"26400000" after 126.5632816408204us,
    X"26400000" after 126.66333166583291us,
    X"26400000" after 126.76338169084542us,
    X"26400000" after 126.86343171585793us,
    X"26400000" after 126.96348174087042us,
    X"26400000" after 127.06353176588293us,
    X"26400000" after 127.16358179089544us,
    X"26400000" after 127.26363181590794us,
    X"26400000" after 127.36368184092045us,
    X"26400000" after 127.46373186593296us,
    X"26400000" after 127.56378189094546us,
    X"26400000" after 127.66383191595797us,
    X"26400000" after 127.76388194097048us,
    X"26400000" after 127.86393196598299us,
    X"26400000" after 127.96398199099549us,
    X"26400000" after 128.06403201600799us,
    X"26400000" after 128.1640820410205us,
    X"26400000" after 128.264132066033us,
    X"26400000" after 128.3641820910455us,
    X"26400000" after 128.464232116058us,
    X"26400000" after 128.56428214107052us,
    X"26400000" after 128.66433216608303us,
    X"26400000" after 128.76438219109554us,
    X"26400000" after 128.86443221610804us,
    X"26400000" after 128.96448224112055us,
    X"26400000" after 129.06453226613306us,
    X"26400000" after 129.16458229114556us,
    X"26400000" after 129.26463231615807us,
    X"26400000" after 129.36468234117058us,
    X"26400000" after 129.46473236618309us,
    X"26400000" after 129.5647823911956us,
    X"26400000" after 129.6648324162081us,
    X"26400000" after 129.7648824412206us,
    X"26400000" after 129.8649324662331us,
    X"26400000" after 129.96498249124562us,
    X"ffffffff" after 130.06503251625813us,
    X"ffffffff" after 130.16508254127064us,
    X"ffffffff" after 130.26513256628314us,
    X"ffffffff" after 130.36518259129565us,
    X"ffffffff" after 130.46523261630816us,
    X"ffffffff" after 130.56528264132066us,
    X"ffffffff" after 130.66533266633317us,
    X"ffffffff" after 130.76538269134568us,
    X"ffffffff" after 130.86543271635816us,
    X"ffffffff" after 130.96548274137066us,
    X"ffffffff" after 131.06553276638317us,
    X"ffffffff" after 131.16558279139568us,
    X"ffffffff" after 131.26563281640819us,
    X"ffffffff" after 131.3656828414207us,
    X"ffffffff" after 131.4657328664332us,
    X"ffffffff" after 131.5657828914457us,
    X"ffffffff" after 131.6658329164582us,
    X"ffffffff" after 131.76588294147072us,
    X"ffffffff" after 131.86593296648323us,
    X"ffffffff" after 131.96598299149574us,
    X"ffffffff" after 132.06603301650824us,
    X"ffffffff" after 132.16608304152075us,
    X"ffffffff" after 132.26613306653326us,
    X"ffffffff" after 132.36618309154576us,
    X"ffffffff" after 132.46623311655827us,
    X"ffffffff" after 132.56628314157078us,
    X"ffffffff" after 132.66633316658329us,
    X"ffffffff" after 132.7663831915958us,
    X"ffffffff" after 132.8664332166083us,
    X"ffffffff" after 132.9664832416208us,
    X"ffffffff" after 133.06653326663331us,
    X"ffffffff" after 133.16658329164582us,
    X"ffffffff" after 133.26663331665833us,
    X"ffffffff" after 133.36668334167084us,
    X"ffffffff" after 133.46673336668334us,
    X"ffffffff" after 133.56678339169585us,
    X"ffffffff" after 133.66683341670836us,
    X"ffffffff" after 133.76688344172086us,
    X"ffffffff" after 133.86693346673337us,
    X"ffffffff" after 133.96698349174588us,
    X"ffffffff" after 134.06703351675836us,
    X"ffffffff" after 134.16708354177086us,
    X"ffffffff" after 134.26713356678337us,
    X"ffffffff" after 134.36718359179588us,
    X"ffffffff" after 134.4672336168084us,
    X"ffffffff" after 134.5672836418209us,
    X"ffffffff" after 134.6673336668334us,
    X"ffffffff" after 134.7673836918459us,
    X"ffffffff" after 134.86743371685841us,
    X"ffffffff" after 134.96748374187092us,
    X"ffffffff" after 135.06753376688343us,
    X"ffffffff" after 135.16758379189594us,
    X"ffffffff" after 135.26763381690844us,
    X"ffffffff" after 135.36768384192095us,
    X"ffffffff" after 135.46773386693346us,
    X"ffffffff" after 135.56778389194596us,
    X"ffffffff" after 135.66783391695847us,
    X"ffffffff" after 135.76788394197098us,
    X"ffffffff" after 135.8679339669835us,
    X"ffffffff" after 135.967983991996us,
    X"ffffffff" after 136.0680340170085us,
    X"ffffffff" after 136.168084042021us,
    X"ffffffff" after 136.26813406703351us,
    X"ffffffff" after 136.36818409204602us,
    X"ffffffff" after 136.46823411705853us,
    X"ffffffff" after 136.56828414207104us,
    X"ffffffff" after 136.66833416708354us,
    X"ffffffff" after 136.76838419209605us,
    X"ffffffff" after 136.86843421710856us,
    X"ffffffff" after 136.96848424212106us,
    X"ffffffff" after 137.06853426713357us,
    X"ffffffff" after 137.16858429214605us,
    X"ffffffff" after 137.26863431715856us,
    X"ffffffff" after 137.36868434217106us,
    X"ffffffff" after 137.46873436718357us,
    X"ffffffff" after 137.56878439219608us,
    X"ffffffff" after 137.6688344172086us,
    X"ffffffff" after 137.7688844422211us,
    X"ffffffff" after 137.8689344672336us,
    X"ffffffff" after 137.9689844922461us,
    X"ffffffff" after 138.06903451725861us,
    X"ffffffff" after 138.16908454227112us,
    X"ffffffff" after 138.26913456728363us,
    X"ffffffff" after 138.36918459229614us,
    X"ffffffff" after 138.46923461730864us,
    X"ffffffff" after 138.56928464232115us,
    X"ffffffff" after 138.66933466733366us,
    X"ffffffff" after 138.76938469234616us,
    X"ffffffff" after 138.86943471735867us,
    X"ffffffff" after 138.96948474237118us,
    X"ffffffff" after 139.0695347673837us,
    X"ffffffff" after 139.1695847923962us,
    X"ffffffff" after 139.2696348174087us,
    X"ffffffff" after 139.3696848424212us,
    X"ffffffff" after 139.46973486743371us,
    X"ffffffff" after 139.56978489244622us,
    X"ffffffff" after 139.66983491745873us,
    X"ffffffff" after 139.76988494247124us,
    X"ffffffff" after 139.86993496748374us,
    X"ffffffff" after 139.96998499249625us,
    X"ffffffff" after 140.07003501750876us,
    X"ffffffff" after 140.17008504252126us,
    X"ffffffff" after 140.27013506753377us,
    X"ffffffff" after 140.37018509254625us,
    X"ffffffff" after 140.47023511755876us,
    X"ffffffff" after 140.57028514257127us,
    X"ffffffff" after 140.67033516758377us,
    X"ffffffff" after 140.77038519259628us,
    X"ffffffff" after 140.8704352176088us,
    X"ffffffff" after 140.9704852426213us,
    X"ffffffff" after 141.0705352676338us,
    X"ffffffff" after 141.1705852926463us,
    X"ffffffff" after 141.27063531765882us,
    X"ffffffff" after 141.37068534267132us,
    X"ffffffff" after 141.47073536768383us,
    X"ffffffff" after 141.57078539269634us,
    X"ffffffff" after 141.67083541770884us,
    X"ffffffff" after 141.77088544272135us,
    X"ffffffff" after 141.87093546773386us,
    X"ffffffff" after 141.97098549274637us,
    X"ffffffff" after 142.07103551775887us,
    X"ffffffff" after 142.17108554277138us,
    X"ffffffff" after 142.2711355677839us,
    X"ffffffff" after 142.3711855927964us,
    X"ffffffff" after 142.4712356178089us,
    X"ffffffff" after 142.5712856428214us,
    X"ffffffff" after 142.67133566783392us,
    X"ffffffff" after 142.77138569284642us,
    X"ffffffff" after 142.87143571785893us,
    X"ffffffff" after 142.97148574287144us,
    X"ffffffff" after 143.07153576788394us,
    X"ffffffff" after 143.17158579289645us,
    X"ffffffff" after 143.27163581790896us,
    X"ffffffff" after 143.37168584292147us,
    X"ffffffff" after 143.47173586793394us,
    X"ffffffff" after 143.57178589294645us,
    X"ffffffff" after 143.67183591795896us,
    X"ffffffff" after 143.77188594297147us,
    X"ffffffff" after 143.87193596798397us,
    X"ffffffff" after 143.97198599299648us,
    X"ffffffff" after 144.072036018009us,
    X"ffffffff" after 144.1720860430215us,
    X"ffffffff" after 144.272136068034us,
    X"ffffffff" after 144.3721860930465us,
    X"ffffffff" after 144.47223611805902us,
    X"ffffffff" after 144.57228614307152us,
    X"ffffffff" after 144.67233616808403us,
    X"ffffffff" after 144.77238619309654us,
    X"ffffffff" after 144.87243621810904us,
    X"ffffffff" after 144.97248624312155us,
    X"ffffffff" after 145.07253626813406us,
    X"ffffffff" after 145.17258629314657us,
    X"ffffffff" after 145.27263631815907us,
    X"ffffffff" after 145.37268634317158us,
    X"ffffffff" after 145.4727363681841us,
    X"ffffffff" after 145.5727863931966us,
    X"ffffffff" after 145.6728364182091us,
    X"ffffffff" after 145.7728864432216us,
    X"ffffffff" after 145.87293646823412us,
    X"ffffffff" after 145.97298649324662us,
    X"ffffffff" after 146.07303651825913us,
    X"ffffffff" after 146.17308654327164us,
    X"ffffffff" after 146.27313656828414us,
    X"ffffffff" after 146.37318659329665us,
    X"ffffffff" after 146.47323661830916us,
    X"ffffffff" after 146.57328664332167us,
    X"ffffffff" after 146.67333666833414us,
    X"ffffffff" after 146.77338669334665us,
    X"ffffffff" after 146.87343671835916us,
    X"ffffffff" after 146.97348674337167us,
    X"ffffffff" after 147.07353676838417us,
    X"ffffffff" after 147.17358679339668us,
    X"ffffffff" after 147.2736368184092us,
    X"ffffffff" after 147.3736868434217us,
    X"ffffffff" after 147.4737368684342us,
    X"ffffffff" after 147.5737868934467us,
    X"ffffffff" after 147.67383691845922us,
    X"ffffffff" after 147.77388694347172us,
    X"ffffffff" after 147.87393696848423us,
    X"ffffffff" after 147.97398699349674us,
    X"ffffffff" after 148.07403701850924us,
    X"ffffffff" after 148.17408704352175us,
    X"ffffffff" after 148.27413706853426us,
    X"ffffffff" after 148.37418709354677us,
    X"ffffffff" after 148.47423711855927us,
    X"ffffffff" after 148.57428714357178us,
    X"ffffffff" after 148.6743371685843us,
    X"ffffffff" after 148.7743871935968us,
    X"ffffffff" after 148.8744372186093us,
    X"ffffffff" after 148.9744872436218us,
    X"ffffffff" after 149.07453726863432us,
    X"ffffffff" after 149.17458729364682us,
    X"ffffffff" after 149.27463731865933us,
    X"ffffffff" after 149.37468734367184us,
    X"ffffffff" after 149.47473736868434us,
    X"ffffffff" after 149.57478739369685us,
    X"ffffffff" after 149.67483741870936us,
    X"ffffffff" after 149.77488744372184us,
    X"ffffffff" after 149.87493746873434us,
    X"ffffffff" after 149.97498749374685us,
    X"80000000" after 150.07503751875936us,
    X"80000000" after 150.17508754377187us,
    X"80000000" after 150.27513756878437us,
    X"80000000" after 150.37518759379688us,
    X"80000000" after 150.4752376188094us,
    X"80000000" after 150.5752876438219us,
    X"80000000" after 150.6753376688344us,
    X"80000000" after 150.7753876938469us,
    X"80000000" after 150.87543771885942us,
    X"80000000" after 150.97548774387192us,
    X"80000000" after 151.07553776888443us,
    X"80000000" after 151.17558779389694us,
    X"80000000" after 151.27563781890944us,
    X"80000000" after 151.37568784392195us,
    X"80000000" after 151.47573786893446us,
    X"80000000" after 151.57578789394697us,
    X"80000000" after 151.67583791895947us,
    X"80000000" after 151.77588794397198us,
    X"80000000" after 151.8759379689845us,
    X"80000000" after 151.975987993997us,
    X"80000000" after 152.0760380190095us,
    X"80000000" after 152.176088044022us,
    X"80000000" after 152.27613806903452us,
    X"80000000" after 152.37618809404702us,
    X"80000000" after 152.47623811905953us,
    X"80000000" after 152.57628814407204us,
    X"80000000" after 152.67633816908454us,
    X"80000000" after 152.77638819409705us,
    X"80000000" after 152.87643821910956us,
    X"80000000" after 152.97648824412204us,
    X"80000000" after 153.07653826913455us,
    X"80000000" after 153.17658829414705us,
    X"80000000" after 153.27663831915956us,
    X"80000000" after 153.37668834417207us,
    X"80000000" after 153.47673836918457us,
    X"80000000" after 153.57678839419708us,
    X"80000000" after 153.6768384192096us,
    X"80000000" after 153.7768884442221us,
    X"80000000" after 153.8769384692346us,
    X"80000000" after 153.9769884942471us,
    X"80000000" after 154.07703851925962us,
    X"80000000" after 154.17708854427212us,
    X"80000000" after 154.27713856928463us,
    X"80000000" after 154.37718859429714us,
    X"80000000" after 154.47723861930965us,
    X"80000000" after 154.57728864432215us,
    X"80000000" after 154.67733866933466us,
    X"80000000" after 154.77738869434717us,
    X"80000000" after 154.87743871935967us,
    X"80000000" after 154.97748874437218us,
    X"80000000" after 155.0775387693847us,
    X"80000000" after 155.1775887943972us,
    X"80000000" after 155.2776388194097us,
    X"80000000" after 155.3776888444222us,
    X"80000000" after 155.47773886943472us,
    X"80000000" after 155.57778889444722us,
    X"80000000" after 155.67783891945973us,
    X"80000000" after 155.77788894447224us,
    X"80000000" after 155.87793896948475us,
    X"80000000" after 155.97798899449725us,
    X"80000000" after 156.07803901950973us,
    X"80000000" after 156.17808904452224us,
    X"80000000" after 156.27813906953475us,
    X"80000000" after 156.37818909454725us,
    X"80000000" after 156.47823911955976us,
    X"80000000" after 156.57828914457227us,
    X"80000000" after 156.67833916958477us,
    X"80000000" after 156.77838919459728us,
    X"80000000" after 156.8784392196098us,
    X"80000000" after 156.9784892446223us,
    X"80000000" after 157.0785392696348us,
    X"80000000" after 157.1785892946473us,
    X"80000000" after 157.27863931965982us,
    X"80000000" after 157.37868934467232us,
    X"80000000" after 157.47873936968483us,
    X"80000000" after 157.57878939469734us,
    X"80000000" after 157.67883941970985us,
    X"80000000" after 157.77888944472235us,
    X"80000000" after 157.87893946973486us,
    X"80000000" after 157.97898949474737us,
    X"80000000" after 158.07903951975987us,
    X"80000000" after 158.17908954477238us,
    X"80000000" after 158.2791395697849us,
    X"80000000" after 158.3791895947974us,
    X"80000000" after 158.4792396198099us,
    X"80000000" after 158.5792896448224us,
    X"80000000" after 158.67933966983492us,
    X"80000000" after 158.77938969484742us,
    X"80000000" after 158.87943971985993us,
    X"80000000" after 158.97948974487244us,
    X"80000000" after 159.07953976988495us,
    X"80000000" after 159.17958979489745us,
    X"80000000" after 159.27963981990993us,
    X"80000000" after 159.37968984492244us,
    X"80000000" after 159.47973986993495us,
    X"80000000" after 159.57978989494745us,
    X"80000000" after 159.67983991995996us,
    X"80000000" after 159.77988994497247us,
    X"80000000" after 159.87993996998497us,
    X"80000000" after 159.97998999499748us,
    X"ffffffff" after 160.08004002001us,
    X"ffffffff" after 160.1800900450225us,
    X"ffffffff" after 160.280140070035us,
    X"ffffffff" after 160.3801900950475us,
    X"ffffffff" after 160.48024012006002us,
    X"ffffffff" after 160.58029014507252us,
    X"ffffffff" after 160.68034017008503us,
    X"ffffffff" after 160.78039019509754us,
    X"ffffffff" after 160.88044022011005us,
    X"ffffffff" after 160.98049024512255us,
    X"ffffffff" after 161.08054027013506us,
    X"ffffffff" after 161.18059029514757us,
    X"ffffffff" after 161.28064032016007us,
    X"ffffffff" after 161.38069034517258us,
    X"ffffffff" after 161.4807403701851us,
    X"ffffffff" after 161.5807903951976us,
    X"ffffffff" after 161.6808404202101us,
    X"ffffffff" after 161.7808904452226us,
    X"ffffffff" after 161.88094047023512us,
    X"ffffffff" after 161.98099049524762us,
    X"ffffffff" after 162.08104052026013us,
    X"ffffffff" after 162.18109054527264us,
    X"ffffffff" after 162.28114057028515us,
    X"ffffffff" after 162.38119059529762us,
    X"ffffffff" after 162.48124062031013us,
    X"ffffffff" after 162.58129064532264us,
    X"ffffffff" after 162.68134067033515us,
    X"ffffffff" after 162.78139069534765us,
    X"ffffffff" after 162.88144072036016us,
    X"ffffffff" after 162.98149074537267us,
    X"ffffffff" after 163.08154077038517us,
    X"ffffffff" after 163.18159079539768us,
    X"ffffffff" after 163.2816408204102us,
    X"ffffffff" after 163.3816908454227us,
    X"ffffffff" after 163.4817408704352us,
    X"ffffffff" after 163.5817908954477us,
    X"ffffffff" after 163.68184092046022us,
    X"ffffffff" after 163.78189094547272us,
    X"ffffffff" after 163.88194097048523us,
    X"ffffffff" after 163.98199099549774us,
    X"ffffffff" after 164.08204102051025us,
    X"ffffffff" after 164.18209104552275us,
    X"ffffffff" after 164.28214107053526us,
    X"ffffffff" after 164.38219109554777us,
    X"ffffffff" after 164.48224112056027us,
    X"ffffffff" after 164.58229114557278us,
    X"ffffffff" after 164.6823411705853us,
    X"ffffffff" after 164.7823911955978us,
    X"ffffffff" after 164.8824412206103us,
    X"ffffffff" after 164.9824912456228us,
    X"ffffffff" after 165.08254127063532us,
    X"ffffffff" after 165.18259129564782us,
    X"ffffffff" after 165.28264132066033us,
    X"ffffffff" after 165.38269134567284us,
    X"ffffffff" after 165.48274137068535us,
    X"ffffffff" after 165.58279139569783us,
    X"ffffffff" after 165.68284142071033us,
    X"ffffffff" after 165.78289144572284us,
    X"ffffffff" after 165.88294147073535us,
    X"ffffffff" after 165.98299149574785us,
    X"ffffffff" after 166.08304152076036us,
    X"ffffffff" after 166.18309154577287us,
    X"ffffffff" after 166.28314157078538us,
    X"ffffffff" after 166.38319159579788us,
    X"ffffffff" after 166.4832416208104us,
    X"ffffffff" after 166.5832916458229us,
    X"ffffffff" after 166.6833416708354us,
    X"ffffffff" after 166.7833916958479us,
    X"ffffffff" after 166.88344172086042us,
    X"ffffffff" after 166.98349174587293us,
    X"ffffffff" after 167.08354177088543us,
    X"ffffffff" after 167.18359179589794us,
    X"ffffffff" after 167.28364182091045us,
    X"ffffffff" after 167.38369184592295us,
    X"ffffffff" after 167.48374187093546us,
    X"ffffffff" after 167.58379189594797us,
    X"ffffffff" after 167.68384192096048us,
    X"ffffffff" after 167.78389194597298us,
    X"ffffffff" after 167.8839419709855us,
    X"ffffffff" after 167.983991995998us,
    X"ffffffff" after 168.0840420210105us,
    X"ffffffff" after 168.184092046023us,
    X"ffffffff" after 168.28414207103552us,
    X"ffffffff" after 168.38419209604803us,
    X"ffffffff" after 168.48424212106053us,
    X"ffffffff" after 168.58429214607304us,
    X"ffffffff" after 168.68434217108552us,
    X"ffffffff" after 168.78439219609803us,
    X"ffffffff" after 168.88444222111053us,
    X"ffffffff" after 168.98449224612304us,
    X"ffffffff" after 169.08454227113555us,
    X"ffffffff" after 169.18459229614805us,
    X"ffffffff" after 169.28464232116056us,
    X"ffffffff" after 169.38469234617307us,
    X"ffffffff" after 169.48474237118558us,
    X"ffffffff" after 169.58479239619808us,
    X"ffffffff" after 169.6848424212106us,
    X"ffffffff" after 169.7848924462231us,
    X"ffffffff" after 169.8849424712356us,
    X"ffffffff" after 169.9849924962481us,
    X"ffffffff" after 170.08504252126062us,
    X"ffffffff" after 170.18509254627313us,
    X"ffffffff" after 170.28514257128563us,
    X"ffffffff" after 170.38519259629814us,
    X"ffffffff" after 170.48524262131065us,
    X"ffffffff" after 170.58529264632315us,
    X"ffffffff" after 170.68534267133566us,
    X"ffffffff" after 170.78539269634817us,
    X"ffffffff" after 170.88544272136068us,
    X"ffffffff" after 170.98549274637318us,
    X"ffffffff" after 171.0855427713857us,
    X"ffffffff" after 171.1855927963982us,
    X"ffffffff" after 171.2856428214107us,
    X"ffffffff" after 171.3856928464232us,
    X"ffffffff" after 171.48574287143572us,
    X"ffffffff" after 171.58579289644823us,
    X"ffffffff" after 171.68584292146073us,
    X"ffffffff" after 171.78589294647324us,
    X"ffffffff" after 171.88594297148572us,
    X"ffffffff" after 171.98599299649823us,
    X"ffffffff" after 172.08604302151073us,
    X"ffffffff" after 172.18609304652324us,
    X"ffffffff" after 172.28614307153575us,
    X"ffffffff" after 172.38619309654825us,
    X"ffffffff" after 172.48624312156076us,
    X"ffffffff" after 172.58629314657327us,
    X"ffffffff" after 172.68634317158578us,
    X"ffffffff" after 172.78639319659828us,
    X"ffffffff" after 172.8864432216108us,
    X"ffffffff" after 172.9864932466233us,
    X"ffffffff" after 173.0865432716358us,
    X"ffffffff" after 173.1865932966483us,
    X"ffffffff" after 173.28664332166082us,
    X"ffffffff" after 173.38669334667333us,
    X"ffffffff" after 173.48674337168583us,
    X"ffffffff" after 173.58679339669834us,
    X"ffffffff" after 173.68684342171085us,
    X"ffffffff" after 173.78689344672335us,
    X"ffffffff" after 173.88694347173586us,
    X"ffffffff" after 173.98699349674837us,
    X"ffffffff" after 174.08704352176088us,
    X"ffffffff" after 174.18709354677338us,
    X"ffffffff" after 174.2871435717859us,
    X"ffffffff" after 174.3871935967984us,
    X"ffffffff" after 174.4872436218109us,
    X"ffffffff" after 174.5872936468234us,
    X"ffffffff" after 174.68734367183592us,
    X"ffffffff" after 174.78739369684843us,
    X"ffffffff" after 174.88744372186093us,
    X"ffffffff" after 174.9874937468734us,
    X"26400000" after 175.08754377188592us,
    X"26400000" after 175.18759379689843us,
    X"26400000" after 175.28764382191093us,
    X"26400000" after 175.38769384692344us,
    X"26400000" after 175.48774387193595us,
    X"26400000" after 175.58779389694845us,
    X"26400000" after 175.68784392196096us,
    X"26400000" after 175.78789394697347us,
    X"26400000" after 175.88794397198598us,
    X"26400000" after 175.98799399699848us,
    X"26400000" after 176.088044022011us,
    X"26400000" after 176.1880940470235us,
    X"26400000" after 176.288144072036us,
    X"26400000" after 176.3881940970485us,
    X"26400000" after 176.48824412206102us,
    X"26400000" after 176.58829414707353us,
    X"26400000" after 176.68834417208603us,
    X"26400000" after 176.78839419709854us,
    X"26400000" after 176.88844422211105us,
    X"26400000" after 176.98849424712355us,
    X"26400000" after 177.08854427213606us,
    X"26400000" after 177.18859429714857us,
    X"26400000" after 177.28864432216108us,
    X"26400000" after 177.38869434717358us,
    X"26400000" after 177.4887443721861us,
    X"26400000" after 177.5887943971986us,
    X"26400000" after 177.6888444222111us,
    X"26400000" after 177.7888944472236us,
    X"26400000" after 177.88894447223612us,
    X"26400000" after 177.98899449724863us,
    X"26400000" after 178.08904452226113us,
    X"26400000" after 178.1890945472736us,
    X"26400000" after 178.28914457228612us,
    X"26400000" after 178.38919459729863us,
    X"26400000" after 178.48924462231113us,
    X"26400000" after 178.58929464732364us,
    X"26400000" after 178.68934467233615us,
    X"26400000" after 178.78939469734865us,
    X"26400000" after 178.88944472236116us,
    X"26400000" after 178.98949474737367us,
    X"26400000" after 179.08954477238618us,
    X"26400000" after 179.18959479739868us,
    X"26400000" after 179.2896448224112us,
    X"26400000" after 179.3896948474237us,
    X"26400000" after 179.4897448724362us,
    X"26400000" after 179.5897948974487us,
    X"26400000" after 179.68984492246122us,
    X"26400000" after 179.78989494747373us,
    X"26400000" after 179.88994497248623us,
    X"26400000" after 179.98999499749874us,
    X"ffffffff" after 180.09004502251125us,
    X"ffffffff" after 180.19009504752376us,
    X"ffffffff" after 180.29014507253626us,
    X"ffffffff" after 180.39019509754877us,
    X"ffffffff" after 180.49024512256128us,
    X"ffffffff" after 180.59029514757378us,
    X"ffffffff" after 180.6903451725863us,
    X"ffffffff" after 180.7903951975988us,
    X"ffffffff" after 180.8904452226113us,
    X"ffffffff" after 180.9904952476238us,
    X"ffffffff" after 181.09054527263632us,
    X"ffffffff" after 181.19059529764883us,
    X"ffffffff" after 181.2906453226613us,
    X"ffffffff" after 181.3906953476738us,
    X"ffffffff" after 181.49074537268632us,
    X"ffffffff" after 181.59079539769883us,
    X"ffffffff" after 181.69084542271133us,
    X"ffffffff" after 181.79089544772384us,
    X"ffffffff" after 181.89094547273635us,
    X"ffffffff" after 181.99099549774886us,
    X"ffffffff" after 182.09104552276136us,
    X"ffffffff" after 182.19109554777387us,
    X"ffffffff" after 182.29114557278638us,
    X"ffffffff" after 182.39119559779888us,
    X"ffffffff" after 182.4912456228114us,
    X"ffffffff" after 182.5912956478239us,
    X"ffffffff" after 182.6913456728364us,
    X"ffffffff" after 182.7913956978489us,
    X"ffffffff" after 182.89144572286142us,
    X"ffffffff" after 182.99149574787393us,
    X"ffffffff" after 183.09154577288643us,
    X"ffffffff" after 183.19159579789894us,
    X"ffffffff" after 183.29164582291145us,
    X"ffffffff" after 183.39169584792396us,
    X"ffffffff" after 183.49174587293646us,
    X"ffffffff" after 183.59179589794897us,
    X"ffffffff" after 183.69184592296148us,
    X"ffffffff" after 183.79189594797398us,
    X"ffffffff" after 183.8919459729865us,
    X"ffffffff" after 183.991995997999us,
    X"ffffffff" after 184.0920460230115us,
    X"ffffffff" after 184.192096048024us,
    X"ffffffff" after 184.29214607303652us,
    X"ffffffff" after 184.39219609804903us,
    X"ffffffff" after 184.4922461230615us,
    X"ffffffff" after 184.592296148074us,
    X"ffffffff" after 184.69234617308652us,
    X"ffffffff" after 184.79239619809903us,
    X"ffffffff" after 184.89244622311153us,
    X"ffffffff" after 184.99249624812404us,
    X"ffffffff" after 185.09254627313655us,
    X"ffffffff" after 185.19259629814906us,
    X"ffffffff" after 185.29264632316156us,
    X"ffffffff" after 185.39269634817407us,
    X"ffffffff" after 185.49274637318658us,
    X"ffffffff" after 185.59279639819908us,
    X"ffffffff" after 185.6928464232116us,
    X"ffffffff" after 185.7928964482241us,
    X"ffffffff" after 185.8929464732366us,
    X"ffffffff" after 185.9929964982491us,
    X"ffffffff" after 186.09304652326162us,
    X"ffffffff" after 186.19309654827413us,
    X"ffffffff" after 186.29314657328663us,
    X"ffffffff" after 186.39319659829914us,
    X"ffffffff" after 186.49324662331165us,
    X"ffffffff" after 186.59329664832416us,
    X"ffffffff" after 186.69334667333666us,
    X"ffffffff" after 186.79339669834917us,
    X"ffffffff" after 186.89344672336168us,
    X"ffffffff" after 186.99349674837418us,
    X"ffffffff" after 187.0935467733867us,
    X"ffffffff" after 187.1935967983992us,
    X"ffffffff" after 187.2936468234117us,
    X"ffffffff" after 187.3936968484242us,
    X"ffffffff" after 187.49374687343672us,
    X"ffffffff" after 187.5937968984492us,
    X"ffffffff" after 187.6938469234617us,
    X"ffffffff" after 187.7938969484742us,
    X"ffffffff" after 187.89394697348672us,
    X"ffffffff" after 187.99399699849923us,
    X"ffffffff" after 188.09404702351173us,
    X"ffffffff" after 188.19409704852424us,
    X"ffffffff" after 188.29414707353675us,
    X"ffffffff" after 188.39419709854926us,
    X"ffffffff" after 188.49424712356176us,
    X"ffffffff" after 188.59429714857427us,
    X"ffffffff" after 188.69434717358678us,
    X"ffffffff" after 188.79439719859928us,
    X"ffffffff" after 188.8944472236118us,
    X"ffffffff" after 188.9944972486243us,
    X"ffffffff" after 189.0945472736368us,
    X"ffffffff" after 189.1945972986493us,
    X"ffffffff" after 189.29464732366182us,
    X"ffffffff" after 189.39469734867433us,
    X"ffffffff" after 189.49474737368683us,
    X"ffffffff" after 189.59479739869934us,
    X"ffffffff" after 189.69484742371185us,
    X"ffffffff" after 189.79489744872436us,
    X"ffffffff" after 189.89494747373686us,
    X"ffffffff" after 189.99499749874937us,
    X"ffffffff" after 190.09504752376188us,
    X"ffffffff" after 190.19509754877438us,
    X"ffffffff" after 190.2951475737869us,
    X"ffffffff" after 190.3951975987994us,
    X"ffffffff" after 190.4952476238119us,
    X"ffffffff" after 190.5952976488244us,
    X"ffffffff" after 190.69534767383692us,
    X"ffffffff" after 190.7953976988494us,
    X"ffffffff" after 190.8954477238619us,
    X"ffffffff" after 190.9954977488744us,
    X"ffffffff" after 191.09554777388692us,
    X"ffffffff" after 191.19559779889943us,
    X"ffffffff" after 191.29564782391193us,
    X"ffffffff" after 191.39569784892444us,
    X"ffffffff" after 191.49574787393695us,
    X"ffffffff" after 191.59579789894946us,
    X"ffffffff" after 191.69584792396196us,
    X"ffffffff" after 191.79589794897447us,
    X"ffffffff" after 191.89594797398698us,
    X"ffffffff" after 191.99599799899948us,
    X"ffffffff" after 192.096048024012us,
    X"ffffffff" after 192.1960980490245us,
    X"ffffffff" after 192.296148074037us,
    X"ffffffff" after 192.3961980990495us,
    X"ffffffff" after 192.49624812406202us,
    X"ffffffff" after 192.59629814907453us,
    X"ffffffff" after 192.69634817408703us,
    X"ffffffff" after 192.79639819909954us,
    X"ffffffff" after 192.89644822411205us,
    X"ffffffff" after 192.99649824912456us,
    X"ffffffff" after 193.09654827413706us,
    X"ffffffff" after 193.19659829914957us,
    X"ffffffff" after 193.29664832416208us,
    X"ffffffff" after 193.39669834917459us,
    X"ffffffff" after 193.4967483741871us,
    X"ffffffff" after 193.5967983991996us,
    X"ffffffff" after 193.6968484242121us,
    X"ffffffff" after 193.7968984492246us,
    X"ffffffff" after 193.8969484742371us,
    X"ffffffff" after 193.9969984992496us,
    X"ffffffff" after 194.0970485242621us,
    X"ffffffff" after 194.1970985492746us,
    X"ffffffff" after 194.29714857428712us,
    X"ffffffff" after 194.39719859929963us,
    X"ffffffff" after 194.49724862431214us,
    X"ffffffff" after 194.59729864932464us,
    X"ffffffff" after 194.69734867433715us,
    X"ffffffff" after 194.79739869934966us,
    X"ffffffff" after 194.89744872436216us,
    X"ffffffff" after 194.99749874937467us,
    X"ffffffff" after 195.09754877438718us,
    X"ffffffff" after 195.19759879939969us,
    X"ffffffff" after 195.2976488244122us,
    X"ffffffff" after 195.3976988494247us,
    X"ffffffff" after 195.4977488744372us,
    X"ffffffff" after 195.5977988994497us,
    X"ffffffff" after 195.69784892446222us,
    X"ffffffff" after 195.79789894947473us,
    X"ffffffff" after 195.89794897448724us,
    X"ffffffff" after 195.99799899949974us,
    X"ffffffff" after 196.09804902451225us,
    X"ffffffff" after 196.19809904952476us,
    X"ffffffff" after 196.29814907453726us,
    X"ffffffff" after 196.39819909954977us,
    X"ffffffff" after 196.49824912456228us,
    X"ffffffff" after 196.59829914957479us,
    X"ffffffff" after 196.6983491745873us,
    X"ffffffff" after 196.7983991995998us,
    X"ffffffff" after 196.8984492246123us,
    X"ffffffff" after 196.9984992496248us,
    X"ffffffff" after 197.0985492746373us,
    X"ffffffff" after 197.1985992996498us,
    X"ffffffff" after 197.2986493246623us,
    X"ffffffff" after 197.3986993496748us,
    X"ffffffff" after 197.49874937468732us,
    X"ffffffff" after 197.59879939969983us,
    X"ffffffff" after 197.69884942471234us,
    X"ffffffff" after 197.79889944972484us,
    X"ffffffff" after 197.89894947473735us,
    X"ffffffff" after 197.99899949974986us,
    X"ffffffff" after 198.09904952476236us,
    X"ffffffff" after 198.19909954977487us,
    X"ffffffff" after 198.29914957478738us,
    X"ffffffff" after 198.39919959979989us,
    X"ffffffff" after 198.4992496248124us,
    X"ffffffff" after 198.5992996498249us,
    X"ffffffff" after 198.6993496748374us,
    X"ffffffff" after 198.79939969984991us,
    X"ffffffff" after 198.89944972486242us,
    X"ffffffff" after 198.99949974987493us,
    X"ffffffff" after 199.09954977488744us,
    X"ffffffff" after 199.19959979989994us,
    X"ffffffff" after 199.29964982491245us,
    X"ffffffff" after 199.39969984992496us,
    X"ffffffff" after 199.49974987493746us,
    X"ffffffff" after 199.59979989994997us,
    X"ffffffff" after 199.69984992496248us,
    X"ffffffff" after 199.79989994997499us,
    X"ffffffff" after 199.8999499749875us,
    X"ffffffff" after 200.0us;*/
  
    
end Behavioral; 
